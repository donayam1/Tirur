`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif

module Memory4( // @[:@3.2]
  input          clock, // @[:@4.4]
  input  [10:0]  io_blockio_addr, // @[:@6.4]
  input  [127:0] io_blockio_wdata, // @[:@6.4]
  input          io_blockio_we, // @[:@6.4]
  input          io_blockio_en, // @[:@6.4]
  output [127:0] io_blockio_rdata, // @[:@6.4]
  output         io_blockio_ready, // @[:@6.4]
  input  [12:0]  io_dataio_addr, // @[:@6.4]
  input  [31:0]  io_dataio_wdata, // @[:@6.4]
  input          io_dataio_we, // @[:@6.4]
  input          io_dataio_en, // @[:@6.4]
  output [31:0]  io_dataio_rdata, // @[:@6.4]
  output         io_dataio_ready // @[:@6.4]
);
  reg [7:0] mem_0 [0:8191]; // @[memory4.scala 14:21:@8.4]
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_61_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_61_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_316_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_316_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_397_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_397_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_478_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_478_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_559_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_559_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_44_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_44_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_44_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_44_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_182_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_182_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_182_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_182_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_216_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_216_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_216_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_216_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_250_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_250_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_250_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_250_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_0__T_284_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_0__T_284_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_284_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_0__T_284_en; // @[memory4.scala 14:21:@8.4]
  wire  _GEN_94;
  reg [12:0] mem_0__T_61_addr_pipe_0;
  reg [31:0] _RAND_1;
  wire  _GEN_96;
  reg [12:0] mem_0__T_316_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [12:0] mem_0__T_397_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [12:0] mem_0__T_478_addr_pipe_0;
  reg [31:0] _RAND_4;
  reg [12:0] mem_0__T_559_addr_pipe_0;
  reg [31:0] _RAND_5;
  wire [12:0] _GEN_110;
  wire [12:0] _GEN_114;
  wire [12:0] _GEN_118;
  wire [12:0] _GEN_122;
  reg [7:0] mem_1 [0:8191]; // @[memory4.scala 14:21:@8.4]
  reg [31:0] _RAND_6;
  wire [7:0] mem_1__T_61_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_61_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_316_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_316_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_397_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_397_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_478_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_478_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_559_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_559_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_44_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_44_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_44_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_44_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_182_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_182_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_182_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_182_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_216_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_216_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_216_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_216_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_250_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_250_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_250_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_250_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_1__T_284_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_1__T_284_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_284_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_1__T_284_en; // @[memory4.scala 14:21:@8.4]
  reg [12:0] mem_1__T_61_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [12:0] mem_1__T_316_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [12:0] mem_1__T_397_addr_pipe_0;
  reg [31:0] _RAND_9;
  reg [12:0] mem_1__T_478_addr_pipe_0;
  reg [31:0] _RAND_10;
  reg [12:0] mem_1__T_559_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] mem_2 [0:8191]; // @[memory4.scala 14:21:@8.4]
  reg [31:0] _RAND_12;
  wire [7:0] mem_2__T_61_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_61_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_316_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_316_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_397_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_397_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_478_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_478_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_559_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_559_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_44_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_44_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_44_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_44_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_182_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_182_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_182_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_182_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_216_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_216_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_216_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_216_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_250_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_250_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_250_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_250_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_2__T_284_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_2__T_284_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_284_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_2__T_284_en; // @[memory4.scala 14:21:@8.4]
  reg [12:0] mem_2__T_61_addr_pipe_0;
  reg [31:0] _RAND_13;
  reg [12:0] mem_2__T_316_addr_pipe_0;
  reg [31:0] _RAND_14;
  reg [12:0] mem_2__T_397_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [12:0] mem_2__T_478_addr_pipe_0;
  reg [31:0] _RAND_16;
  reg [12:0] mem_2__T_559_addr_pipe_0;
  reg [31:0] _RAND_17;
  reg [7:0] mem_3 [0:8191]; // @[memory4.scala 14:21:@8.4]
  reg [31:0] _RAND_18;
  wire [7:0] mem_3__T_61_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_61_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_316_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_316_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_397_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_397_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_478_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_478_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_559_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_559_addr; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_44_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_44_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_44_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_44_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_182_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_182_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_182_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_182_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_216_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_216_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_216_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_216_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_250_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_250_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_250_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_250_en; // @[memory4.scala 14:21:@8.4]
  wire [7:0] mem_3__T_284_data; // @[memory4.scala 14:21:@8.4]
  wire [12:0] mem_3__T_284_addr; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_284_mask; // @[memory4.scala 14:21:@8.4]
  wire  mem_3__T_284_en; // @[memory4.scala 14:21:@8.4]
  reg [12:0] mem_3__T_61_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [12:0] mem_3__T_316_addr_pipe_0;
  reg [31:0] _RAND_20;
  reg [12:0] mem_3__T_397_addr_pipe_0;
  reg [31:0] _RAND_21;
  reg [12:0] mem_3__T_478_addr_pipe_0;
  reg [31:0] _RAND_22;
  reg [12:0] mem_3__T_559_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg  _T_74; // @[package.scala 15:91:@44.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_92_0; // @[Reg.scala 11:16:@46.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_92_1; // @[Reg.scala 11:16:@46.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_92_2; // @[Reg.scala 11:16:@46.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_92_3; // @[Reg.scala 11:16:@46.4]
  reg [31:0] _RAND_28;
  reg  _T_329; // @[package.scala 15:91:@203.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_347_0; // @[Reg.scala 11:16:@205.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_347_1; // @[Reg.scala 11:16:@205.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_347_2; // @[Reg.scala 11:16:@205.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_347_3; // @[Reg.scala 11:16:@205.4]
  reg [31:0] _RAND_33;
  reg  _T_410; // @[package.scala 15:91:@228.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_428_0; // @[Reg.scala 11:16:@230.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_428_1; // @[Reg.scala 11:16:@230.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_428_2; // @[Reg.scala 11:16:@230.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_428_3; // @[Reg.scala 11:16:@230.4]
  reg [31:0] _RAND_38;
  reg  _T_491; // @[package.scala 15:91:@253.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_509_0; // @[Reg.scala 11:16:@255.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_509_1; // @[Reg.scala 11:16:@255.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_509_2; // @[Reg.scala 11:16:@255.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_509_3; // @[Reg.scala 11:16:@255.4]
  reg [31:0] _RAND_43;
  reg  _T_572; // @[package.scala 15:91:@278.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_590_0; // @[Reg.scala 11:16:@280.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_590_1; // @[Reg.scala 11:16:@280.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_590_2; // @[Reg.scala 11:16:@280.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_590_3; // @[Reg.scala 11:16:@280.4]
  reg [31:0] _RAND_48;
  wire  wend; // @[memory4.scala 17:29:@9.4]
  wire  _T_27; // @[memory4.scala 18:32:@10.4]
  wire  rend; // @[memory4.scala 18:29:@11.4]
  wire [7:0] datad_0; // @[memory4.scala 22:55:@12.4]
  wire [7:0] datad_1; // @[memory4.scala 22:55:@13.4]
  wire [7:0] datad_2; // @[memory4.scala 22:55:@14.4]
  wire [7:0] datad_3; // @[memory4.scala 22:55:@15.4]
  wire [7:0] _GEN_17; // @[Reg.scala 12:19:@47.4]
  wire [7:0] _GEN_18; // @[Reg.scala 12:19:@47.4]
  wire [7:0] _GEN_19; // @[Reg.scala 12:19:@47.4]
  wire [7:0] _GEN_20; // @[Reg.scala 12:19:@47.4]
  wire [15:0] _T_130; // @[memory4.scala 29:27:@54.4]
  wire [15:0] _T_131; // @[memory4.scala 29:27:@55.4]
  wire [31:0] _T_132; // @[memory4.scala 29:27:@56.4]
  wire  wenb; // @[memory4.scala 37:30:@59.4]
  wire  _T_134; // @[memory4.scala 38:33:@60.4]
  wire  renb; // @[memory4.scala 38:30:@61.4]
  wire [12:0] baseAddr; // @[Cat.scala 30:58:@62.4]
  wire [13:0] _T_161; // @[memory4.scala 52:30:@74.6]
  wire [31:0] _T_163; // @[memory4.scala 53:38:@77.6]
  wire  _T_164; // @[memory4.scala 54:24:@79.6]
  wire [31:0] datab_0; // @[memory4.scala 48:5:@73.4]
  wire [7:0] _T_165; // @[memory4.scala 54:60:@80.6]
  wire [7:0] _T_166; // @[memory4.scala 54:60:@81.6]
  wire [7:0] _T_167; // @[memory4.scala 54:60:@82.6]
  wire [7:0] _T_168; // @[memory4.scala 54:60:@83.6]
  wire [13:0] _T_195; // @[memory4.scala 52:30:@102.6]
  wire [31:0] _T_197; // @[memory4.scala 53:38:@105.6]
  wire  _T_198; // @[memory4.scala 54:24:@107.6]
  wire [31:0] datab_1; // @[memory4.scala 48:5:@73.4]
  wire [7:0] _T_199; // @[memory4.scala 54:60:@108.6]
  wire [7:0] _T_200; // @[memory4.scala 54:60:@109.6]
  wire [7:0] _T_201; // @[memory4.scala 54:60:@110.6]
  wire [7:0] _T_202; // @[memory4.scala 54:60:@111.6]
  wire [13:0] _T_229; // @[memory4.scala 52:30:@130.6]
  wire [31:0] _T_231; // @[memory4.scala 53:38:@133.6]
  wire  _T_232; // @[memory4.scala 54:24:@135.6]
  wire [31:0] datab_2; // @[memory4.scala 48:5:@73.4]
  wire [7:0] _T_233; // @[memory4.scala 54:60:@136.6]
  wire [7:0] _T_234; // @[memory4.scala 54:60:@137.6]
  wire [7:0] _T_235; // @[memory4.scala 54:60:@138.6]
  wire [7:0] _T_236; // @[memory4.scala 54:60:@139.6]
  wire [13:0] _T_263; // @[memory4.scala 52:30:@158.6]
  wire [31:0] _T_265; // @[memory4.scala 53:38:@161.6]
  wire  _T_266; // @[memory4.scala 54:24:@163.6]
  wire [31:0] datab_3; // @[memory4.scala 48:5:@73.4]
  wire [7:0] _T_267; // @[memory4.scala 54:60:@164.6]
  wire [7:0] _T_268; // @[memory4.scala 54:60:@165.6]
  wire [7:0] _T_269; // @[memory4.scala 54:60:@166.6]
  wire [7:0] _T_270; // @[memory4.scala 54:60:@167.6]
  wire [12:0] addrb_0; // @[memory4.scala 63:30:@193.4]
  wire [7:0] _GEN_72; // @[Reg.scala 12:19:@206.4]
  wire [7:0] _GEN_73; // @[Reg.scala 12:19:@206.4]
  wire [7:0] _GEN_74; // @[Reg.scala 12:19:@206.4]
  wire [7:0] _GEN_75; // @[Reg.scala 12:19:@206.4]
  wire [15:0] _T_386; // @[memory4.scala 64:50:@213.4]
  wire [15:0] _T_387; // @[memory4.scala 64:50:@214.4]
  wire [31:0] out_0; // @[memory4.scala 64:50:@215.4]
  wire [12:0] addrb_1; // @[memory4.scala 63:30:@218.4]
  wire [7:0] _GEN_78; // @[Reg.scala 12:19:@231.4]
  wire [7:0] _GEN_79; // @[Reg.scala 12:19:@231.4]
  wire [7:0] _GEN_80; // @[Reg.scala 12:19:@231.4]
  wire [7:0] _GEN_81; // @[Reg.scala 12:19:@231.4]
  wire [15:0] _T_467; // @[memory4.scala 64:50:@238.4]
  wire [15:0] _T_468; // @[memory4.scala 64:50:@239.4]
  wire [31:0] out_1; // @[memory4.scala 64:50:@240.4]
  wire [12:0] addrb_2; // @[memory4.scala 63:30:@243.4]
  wire [7:0] _GEN_84; // @[Reg.scala 12:19:@256.4]
  wire [7:0] _GEN_85; // @[Reg.scala 12:19:@256.4]
  wire [7:0] _GEN_86; // @[Reg.scala 12:19:@256.4]
  wire [7:0] _GEN_87; // @[Reg.scala 12:19:@256.4]
  wire [15:0] _T_548; // @[memory4.scala 64:50:@263.4]
  wire [15:0] _T_549; // @[memory4.scala 64:50:@264.4]
  wire [31:0] out_2; // @[memory4.scala 64:50:@265.4]
  wire [12:0] addrb_3; // @[memory4.scala 63:30:@268.4]
  wire [7:0] _GEN_90; // @[Reg.scala 12:19:@281.4]
  wire [7:0] _GEN_91; // @[Reg.scala 12:19:@281.4]
  wire [7:0] _GEN_92; // @[Reg.scala 12:19:@281.4]
  wire [7:0] _GEN_93; // @[Reg.scala 12:19:@281.4]
  wire [15:0] _T_629; // @[memory4.scala 64:50:@288.4]
  wire [15:0] _T_630; // @[memory4.scala 64:50:@289.4]
  wire [31:0] out_3; // @[memory4.scala 64:50:@290.4]
  wire [63:0] _T_632; // @[Cat.scala 30:58:@292.4]
  wire [63:0] _T_633; // @[Cat.scala 30:58:@293.4]
  wire [127:0] _T_634; // @[Cat.scala 30:58:@294.4]
  assign mem_0__T_61_addr = mem_0__T_61_addr_pipe_0;
  assign mem_0__T_61_data = mem_0[mem_0__T_61_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_0__T_316_addr = mem_0__T_316_addr_pipe_0;
  assign mem_0__T_316_data = mem_0[mem_0__T_316_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_0__T_397_addr = mem_0__T_397_addr_pipe_0;
  assign mem_0__T_397_data = mem_0[mem_0__T_397_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_0__T_478_addr = mem_0__T_478_addr_pipe_0;
  assign mem_0__T_478_data = mem_0[mem_0__T_478_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_0__T_559_addr = mem_0__T_559_addr_pipe_0;
  assign mem_0__T_559_data = mem_0[mem_0__T_559_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_0__T_44_data = datad_0;
  assign mem_0__T_44_addr = io_dataio_addr;
  assign mem_0__T_44_mask = wend;
  assign mem_0__T_44_en = wend;
  assign mem_0__T_182_data = _T_165;
  assign mem_0__T_182_addr = _GEN_110;
  assign mem_0__T_182_mask = wenb;
  assign mem_0__T_182_en = wenb;
  assign mem_0__T_216_data = _T_199;
  assign mem_0__T_216_addr = _GEN_114;
  assign mem_0__T_216_mask = wenb;
  assign mem_0__T_216_en = wenb;
  assign mem_0__T_250_data = _T_233;
  assign mem_0__T_250_addr = _GEN_118;
  assign mem_0__T_250_mask = wenb;
  assign mem_0__T_250_en = wenb;
  assign mem_0__T_284_data = _T_267;
  assign mem_0__T_284_addr = _GEN_122;
  assign mem_0__T_284_mask = wenb;
  assign mem_0__T_284_en = wenb;
  assign _GEN_94 = rend;
  assign _GEN_96 = renb;
  assign _GEN_110 = {{12'd0}, _T_164};
  assign _GEN_114 = {{12'd0}, _T_198};
  assign _GEN_118 = {{12'd0}, _T_232};
  assign _GEN_122 = {{12'd0}, _T_266};
  assign mem_1__T_61_addr = mem_1__T_61_addr_pipe_0;
  assign mem_1__T_61_data = mem_1[mem_1__T_61_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_1__T_316_addr = mem_1__T_316_addr_pipe_0;
  assign mem_1__T_316_data = mem_1[mem_1__T_316_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_1__T_397_addr = mem_1__T_397_addr_pipe_0;
  assign mem_1__T_397_data = mem_1[mem_1__T_397_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_1__T_478_addr = mem_1__T_478_addr_pipe_0;
  assign mem_1__T_478_data = mem_1[mem_1__T_478_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_1__T_559_addr = mem_1__T_559_addr_pipe_0;
  assign mem_1__T_559_data = mem_1[mem_1__T_559_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_1__T_44_data = datad_1;
  assign mem_1__T_44_addr = io_dataio_addr;
  assign mem_1__T_44_mask = wend;
  assign mem_1__T_44_en = wend;
  assign mem_1__T_182_data = _T_166;
  assign mem_1__T_182_addr = _GEN_110;
  assign mem_1__T_182_mask = wenb;
  assign mem_1__T_182_en = wenb;
  assign mem_1__T_216_data = _T_200;
  assign mem_1__T_216_addr = _GEN_114;
  assign mem_1__T_216_mask = wenb;
  assign mem_1__T_216_en = wenb;
  assign mem_1__T_250_data = _T_234;
  assign mem_1__T_250_addr = _GEN_118;
  assign mem_1__T_250_mask = wenb;
  assign mem_1__T_250_en = wenb;
  assign mem_1__T_284_data = _T_268;
  assign mem_1__T_284_addr = _GEN_122;
  assign mem_1__T_284_mask = wenb;
  assign mem_1__T_284_en = wenb;
  assign mem_2__T_61_addr = mem_2__T_61_addr_pipe_0;
  assign mem_2__T_61_data = mem_2[mem_2__T_61_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_2__T_316_addr = mem_2__T_316_addr_pipe_0;
  assign mem_2__T_316_data = mem_2[mem_2__T_316_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_2__T_397_addr = mem_2__T_397_addr_pipe_0;
  assign mem_2__T_397_data = mem_2[mem_2__T_397_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_2__T_478_addr = mem_2__T_478_addr_pipe_0;
  assign mem_2__T_478_data = mem_2[mem_2__T_478_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_2__T_559_addr = mem_2__T_559_addr_pipe_0;
  assign mem_2__T_559_data = mem_2[mem_2__T_559_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_2__T_44_data = datad_2;
  assign mem_2__T_44_addr = io_dataio_addr;
  assign mem_2__T_44_mask = wend;
  assign mem_2__T_44_en = wend;
  assign mem_2__T_182_data = _T_167;
  assign mem_2__T_182_addr = _GEN_110;
  assign mem_2__T_182_mask = wenb;
  assign mem_2__T_182_en = wenb;
  assign mem_2__T_216_data = _T_201;
  assign mem_2__T_216_addr = _GEN_114;
  assign mem_2__T_216_mask = wenb;
  assign mem_2__T_216_en = wenb;
  assign mem_2__T_250_data = _T_235;
  assign mem_2__T_250_addr = _GEN_118;
  assign mem_2__T_250_mask = wenb;
  assign mem_2__T_250_en = wenb;
  assign mem_2__T_284_data = _T_269;
  assign mem_2__T_284_addr = _GEN_122;
  assign mem_2__T_284_mask = wenb;
  assign mem_2__T_284_en = wenb;
  assign mem_3__T_61_addr = mem_3__T_61_addr_pipe_0;
  assign mem_3__T_61_data = mem_3[mem_3__T_61_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_3__T_316_addr = mem_3__T_316_addr_pipe_0;
  assign mem_3__T_316_data = mem_3[mem_3__T_316_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_3__T_397_addr = mem_3__T_397_addr_pipe_0;
  assign mem_3__T_397_data = mem_3[mem_3__T_397_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_3__T_478_addr = mem_3__T_478_addr_pipe_0;
  assign mem_3__T_478_data = mem_3[mem_3__T_478_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_3__T_559_addr = mem_3__T_559_addr_pipe_0;
  assign mem_3__T_559_data = mem_3[mem_3__T_559_addr]; // @[memory4.scala 14:21:@8.4]
  assign mem_3__T_44_data = datad_3;
  assign mem_3__T_44_addr = io_dataio_addr;
  assign mem_3__T_44_mask = wend;
  assign mem_3__T_44_en = wend;
  assign mem_3__T_182_data = _T_168;
  assign mem_3__T_182_addr = _GEN_110;
  assign mem_3__T_182_mask = wenb;
  assign mem_3__T_182_en = wenb;
  assign mem_3__T_216_data = _T_202;
  assign mem_3__T_216_addr = _GEN_114;
  assign mem_3__T_216_mask = wenb;
  assign mem_3__T_216_en = wenb;
  assign mem_3__T_250_data = _T_236;
  assign mem_3__T_250_addr = _GEN_118;
  assign mem_3__T_250_mask = wenb;
  assign mem_3__T_250_en = wenb;
  assign mem_3__T_284_data = _T_270;
  assign mem_3__T_284_addr = _GEN_122;
  assign mem_3__T_284_mask = wenb;
  assign mem_3__T_284_en = wenb;
  assign wend = io_dataio_en & io_dataio_we; // @[memory4.scala 17:29:@9.4]
  assign _T_27 = io_dataio_we == 1'h0; // @[memory4.scala 18:32:@10.4]
  assign rend = io_dataio_en & _T_27; // @[memory4.scala 18:29:@11.4]
  assign datad_0 = io_dataio_wdata[7:0]; // @[memory4.scala 22:55:@12.4]
  assign datad_1 = io_dataio_wdata[15:8]; // @[memory4.scala 22:55:@13.4]
  assign datad_2 = io_dataio_wdata[23:16]; // @[memory4.scala 22:55:@14.4]
  assign datad_3 = io_dataio_wdata[31:24]; // @[memory4.scala 22:55:@15.4]
  assign _GEN_17 = _T_74 ? mem_0__T_61_data : _T_92_0; // @[Reg.scala 12:19:@47.4]
  assign _GEN_18 = _T_74 ? mem_1__T_61_data : _T_92_1; // @[Reg.scala 12:19:@47.4]
  assign _GEN_19 = _T_74 ? mem_2__T_61_data : _T_92_2; // @[Reg.scala 12:19:@47.4]
  assign _GEN_20 = _T_74 ? mem_3__T_61_data : _T_92_3; // @[Reg.scala 12:19:@47.4]
  assign _T_130 = {_GEN_18,_GEN_17}; // @[memory4.scala 29:27:@54.4]
  assign _T_131 = {_GEN_20,_GEN_19}; // @[memory4.scala 29:27:@55.4]
  assign _T_132 = {_T_131,_T_130}; // @[memory4.scala 29:27:@56.4]
  assign wenb = io_blockio_en & io_blockio_we; // @[memory4.scala 37:30:@59.4]
  assign _T_134 = io_blockio_we == 1'h0; // @[memory4.scala 38:33:@60.4]
  assign renb = io_blockio_en & _T_134; // @[memory4.scala 38:30:@61.4]
  assign baseAddr = {io_blockio_addr,2'h0}; // @[Cat.scala 30:58:@62.4]
  assign _T_161 = baseAddr + 13'h0; // @[memory4.scala 52:30:@74.6]
  assign _T_163 = io_blockio_wdata[31:0]; // @[memory4.scala 53:38:@77.6]
  assign _T_164 = io_dataio_addr[0]; // @[memory4.scala 54:24:@79.6]
  assign datab_0 = wenb ? _T_163 : 32'h0; // @[memory4.scala 48:5:@73.4]
  assign _T_165 = datab_0[7:0]; // @[memory4.scala 54:60:@80.6]
  assign _T_166 = datab_0[15:8]; // @[memory4.scala 54:60:@81.6]
  assign _T_167 = datab_0[23:16]; // @[memory4.scala 54:60:@82.6]
  assign _T_168 = datab_0[31:24]; // @[memory4.scala 54:60:@83.6]
  assign _T_195 = baseAddr + 13'h1; // @[memory4.scala 52:30:@102.6]
  assign _T_197 = io_blockio_wdata[63:32]; // @[memory4.scala 53:38:@105.6]
  assign _T_198 = io_dataio_addr[1]; // @[memory4.scala 54:24:@107.6]
  assign datab_1 = wenb ? _T_197 : 32'h0; // @[memory4.scala 48:5:@73.4]
  assign _T_199 = datab_1[7:0]; // @[memory4.scala 54:60:@108.6]
  assign _T_200 = datab_1[15:8]; // @[memory4.scala 54:60:@109.6]
  assign _T_201 = datab_1[23:16]; // @[memory4.scala 54:60:@110.6]
  assign _T_202 = datab_1[31:24]; // @[memory4.scala 54:60:@111.6]
  assign _T_229 = baseAddr + 13'h2; // @[memory4.scala 52:30:@130.6]
  assign _T_231 = io_blockio_wdata[95:64]; // @[memory4.scala 53:38:@133.6]
  assign _T_232 = io_dataio_addr[2]; // @[memory4.scala 54:24:@135.6]
  assign datab_2 = wenb ? _T_231 : 32'h0; // @[memory4.scala 48:5:@73.4]
  assign _T_233 = datab_2[7:0]; // @[memory4.scala 54:60:@136.6]
  assign _T_234 = datab_2[15:8]; // @[memory4.scala 54:60:@137.6]
  assign _T_235 = datab_2[23:16]; // @[memory4.scala 54:60:@138.6]
  assign _T_236 = datab_2[31:24]; // @[memory4.scala 54:60:@139.6]
  assign _T_263 = baseAddr + 13'h3; // @[memory4.scala 52:30:@158.6]
  assign _T_265 = io_blockio_wdata[127:96]; // @[memory4.scala 53:38:@161.6]
  assign _T_266 = io_dataio_addr[3]; // @[memory4.scala 54:24:@163.6]
  assign datab_3 = wenb ? _T_265 : 32'h0; // @[memory4.scala 48:5:@73.4]
  assign _T_267 = datab_3[7:0]; // @[memory4.scala 54:60:@164.6]
  assign _T_268 = datab_3[15:8]; // @[memory4.scala 54:60:@165.6]
  assign _T_269 = datab_3[23:16]; // @[memory4.scala 54:60:@166.6]
  assign _T_270 = datab_3[31:24]; // @[memory4.scala 54:60:@167.6]
  assign addrb_0 = _T_161[12:0]; // @[memory4.scala 63:30:@193.4]
  assign _GEN_72 = _T_329 ? mem_0__T_316_data : _T_347_0; // @[Reg.scala 12:19:@206.4]
  assign _GEN_73 = _T_329 ? mem_1__T_316_data : _T_347_1; // @[Reg.scala 12:19:@206.4]
  assign _GEN_74 = _T_329 ? mem_2__T_316_data : _T_347_2; // @[Reg.scala 12:19:@206.4]
  assign _GEN_75 = _T_329 ? mem_3__T_316_data : _T_347_3; // @[Reg.scala 12:19:@206.4]
  assign _T_386 = {_GEN_73,_GEN_72}; // @[memory4.scala 64:50:@213.4]
  assign _T_387 = {_GEN_75,_GEN_74}; // @[memory4.scala 64:50:@214.4]
  assign out_0 = {_T_387,_T_386}; // @[memory4.scala 64:50:@215.4]
  assign addrb_1 = _T_195[12:0]; // @[memory4.scala 63:30:@218.4]
  assign _GEN_78 = _T_410 ? mem_0__T_397_data : _T_428_0; // @[Reg.scala 12:19:@231.4]
  assign _GEN_79 = _T_410 ? mem_1__T_397_data : _T_428_1; // @[Reg.scala 12:19:@231.4]
  assign _GEN_80 = _T_410 ? mem_2__T_397_data : _T_428_2; // @[Reg.scala 12:19:@231.4]
  assign _GEN_81 = _T_410 ? mem_3__T_397_data : _T_428_3; // @[Reg.scala 12:19:@231.4]
  assign _T_467 = {_GEN_79,_GEN_78}; // @[memory4.scala 64:50:@238.4]
  assign _T_468 = {_GEN_81,_GEN_80}; // @[memory4.scala 64:50:@239.4]
  assign out_1 = {_T_468,_T_467}; // @[memory4.scala 64:50:@240.4]
  assign addrb_2 = _T_229[12:0]; // @[memory4.scala 63:30:@243.4]
  assign _GEN_84 = _T_491 ? mem_0__T_478_data : _T_509_0; // @[Reg.scala 12:19:@256.4]
  assign _GEN_85 = _T_491 ? mem_1__T_478_data : _T_509_1; // @[Reg.scala 12:19:@256.4]
  assign _GEN_86 = _T_491 ? mem_2__T_478_data : _T_509_2; // @[Reg.scala 12:19:@256.4]
  assign _GEN_87 = _T_491 ? mem_3__T_478_data : _T_509_3; // @[Reg.scala 12:19:@256.4]
  assign _T_548 = {_GEN_85,_GEN_84}; // @[memory4.scala 64:50:@263.4]
  assign _T_549 = {_GEN_87,_GEN_86}; // @[memory4.scala 64:50:@264.4]
  assign out_2 = {_T_549,_T_548}; // @[memory4.scala 64:50:@265.4]
  assign addrb_3 = _T_263[12:0]; // @[memory4.scala 63:30:@268.4]
  assign _GEN_90 = _T_572 ? mem_0__T_559_data : _T_590_0; // @[Reg.scala 12:19:@281.4]
  assign _GEN_91 = _T_572 ? mem_1__T_559_data : _T_590_1; // @[Reg.scala 12:19:@281.4]
  assign _GEN_92 = _T_572 ? mem_2__T_559_data : _T_590_2; // @[Reg.scala 12:19:@281.4]
  assign _GEN_93 = _T_572 ? mem_3__T_559_data : _T_590_3; // @[Reg.scala 12:19:@281.4]
  assign _T_629 = {_GEN_91,_GEN_90}; // @[memory4.scala 64:50:@288.4]
  assign _T_630 = {_GEN_93,_GEN_92}; // @[memory4.scala 64:50:@289.4]
  assign out_3 = {_T_630,_T_629}; // @[memory4.scala 64:50:@290.4]
  assign _T_632 = {out_1,out_0}; // @[Cat.scala 30:58:@292.4]
  assign _T_633 = {out_3,out_2}; // @[Cat.scala 30:58:@293.4]
  assign _T_634 = {_T_633,_T_632}; // @[Cat.scala 30:58:@294.4]
  assign io_blockio_rdata = _T_634;
  assign io_blockio_ready = io_blockio_en;
  assign io_dataio_rdata = _T_132;
  assign io_dataio_ready = io_dataio_en;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  _RAND_0 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  mem_0__T_61_addr_pipe_0 = _RAND_1[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  mem_0__T_316_addr_pipe_0 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  mem_0__T_397_addr_pipe_0 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  mem_0__T_478_addr_pipe_0 = _RAND_4[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  mem_0__T_559_addr_pipe_0 = _RAND_5[12:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    mem_1[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  mem_1__T_61_addr_pipe_0 = _RAND_7[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  mem_1__T_316_addr_pipe_0 = _RAND_8[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  mem_1__T_397_addr_pipe_0 = _RAND_9[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  mem_1__T_478_addr_pipe_0 = _RAND_10[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  mem_1__T_559_addr_pipe_0 = _RAND_11[12:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    mem_2[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  mem_2__T_61_addr_pipe_0 = _RAND_13[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  mem_2__T_316_addr_pipe_0 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  mem_2__T_397_addr_pipe_0 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  mem_2__T_478_addr_pipe_0 = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  mem_2__T_559_addr_pipe_0 = _RAND_17[12:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    mem_3[initvar] = _RAND_18[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  mem_3__T_61_addr_pipe_0 = _RAND_19[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  mem_3__T_316_addr_pipe_0 = _RAND_20[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  mem_3__T_397_addr_pipe_0 = _RAND_21[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  mem_3__T_478_addr_pipe_0 = _RAND_22[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  mem_3__T_559_addr_pipe_0 = _RAND_23[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_74 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_92_0 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_92_1 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_92_2 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_92_3 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_329 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_347_0 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_347_1 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_347_2 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_347_3 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_410 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_428_0 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_428_1 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_428_2 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_428_3 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_491 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_509_0 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_509_1 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_509_2 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_509_3 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_572 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_590_0 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_590_1 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_590_2 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_590_3 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem_0__T_44_en & mem_0__T_44_mask) begin
      mem_0[mem_0__T_44_addr] <= mem_0__T_44_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_0__T_182_en & mem_0__T_182_mask) begin
      mem_0[mem_0__T_182_addr] <= mem_0__T_182_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_0__T_216_en & mem_0__T_216_mask) begin
      mem_0[mem_0__T_216_addr] <= mem_0__T_216_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_0__T_250_en & mem_0__T_250_mask) begin
      mem_0[mem_0__T_250_addr] <= mem_0__T_250_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_0__T_284_en & mem_0__T_284_mask) begin
      mem_0[mem_0__T_284_addr] <= mem_0__T_284_data; // @[memory4.scala 14:21:@8.4]
    end
    if (_GEN_94) begin
      mem_0__T_61_addr_pipe_0 <= io_dataio_addr;
    end
    if (_GEN_96) begin
      mem_0__T_316_addr_pipe_0 <= addrb_0;
    end
    if (_GEN_96) begin
      mem_0__T_397_addr_pipe_0 <= addrb_1;
    end
    if (_GEN_96) begin
      mem_0__T_478_addr_pipe_0 <= addrb_2;
    end
    if (_GEN_96) begin
      mem_0__T_559_addr_pipe_0 <= addrb_3;
    end
    if(mem_1__T_44_en & mem_1__T_44_mask) begin
      mem_1[mem_1__T_44_addr] <= mem_1__T_44_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_1__T_182_en & mem_1__T_182_mask) begin
      mem_1[mem_1__T_182_addr] <= mem_1__T_182_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_1__T_216_en & mem_1__T_216_mask) begin
      mem_1[mem_1__T_216_addr] <= mem_1__T_216_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_1__T_250_en & mem_1__T_250_mask) begin
      mem_1[mem_1__T_250_addr] <= mem_1__T_250_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_1__T_284_en & mem_1__T_284_mask) begin
      mem_1[mem_1__T_284_addr] <= mem_1__T_284_data; // @[memory4.scala 14:21:@8.4]
    end
    if (_GEN_94) begin
      mem_1__T_61_addr_pipe_0 <= io_dataio_addr;
    end
    if (_GEN_96) begin
      mem_1__T_316_addr_pipe_0 <= addrb_0;
    end
    if (_GEN_96) begin
      mem_1__T_397_addr_pipe_0 <= addrb_1;
    end
    if (_GEN_96) begin
      mem_1__T_478_addr_pipe_0 <= addrb_2;
    end
    if (_GEN_96) begin
      mem_1__T_559_addr_pipe_0 <= addrb_3;
    end
    if(mem_2__T_44_en & mem_2__T_44_mask) begin
      mem_2[mem_2__T_44_addr] <= mem_2__T_44_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_2__T_182_en & mem_2__T_182_mask) begin
      mem_2[mem_2__T_182_addr] <= mem_2__T_182_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_2__T_216_en & mem_2__T_216_mask) begin
      mem_2[mem_2__T_216_addr] <= mem_2__T_216_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_2__T_250_en & mem_2__T_250_mask) begin
      mem_2[mem_2__T_250_addr] <= mem_2__T_250_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_2__T_284_en & mem_2__T_284_mask) begin
      mem_2[mem_2__T_284_addr] <= mem_2__T_284_data; // @[memory4.scala 14:21:@8.4]
    end
    if (_GEN_94) begin
      mem_2__T_61_addr_pipe_0 <= io_dataio_addr;
    end
    if (_GEN_96) begin
      mem_2__T_316_addr_pipe_0 <= addrb_0;
    end
    if (_GEN_96) begin
      mem_2__T_397_addr_pipe_0 <= addrb_1;
    end
    if (_GEN_96) begin
      mem_2__T_478_addr_pipe_0 <= addrb_2;
    end
    if (_GEN_96) begin
      mem_2__T_559_addr_pipe_0 <= addrb_3;
    end
    if(mem_3__T_44_en & mem_3__T_44_mask) begin
      mem_3[mem_3__T_44_addr] <= mem_3__T_44_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_3__T_182_en & mem_3__T_182_mask) begin
      mem_3[mem_3__T_182_addr] <= mem_3__T_182_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_3__T_216_en & mem_3__T_216_mask) begin
      mem_3[mem_3__T_216_addr] <= mem_3__T_216_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_3__T_250_en & mem_3__T_250_mask) begin
      mem_3[mem_3__T_250_addr] <= mem_3__T_250_data; // @[memory4.scala 14:21:@8.4]
    end
    if(mem_3__T_284_en & mem_3__T_284_mask) begin
      mem_3[mem_3__T_284_addr] <= mem_3__T_284_data; // @[memory4.scala 14:21:@8.4]
    end
    if (_GEN_94) begin
      mem_3__T_61_addr_pipe_0 <= io_dataio_addr;
    end
    if (_GEN_96) begin
      mem_3__T_316_addr_pipe_0 <= addrb_0;
    end
    if (_GEN_96) begin
      mem_3__T_397_addr_pipe_0 <= addrb_1;
    end
    if (_GEN_96) begin
      mem_3__T_478_addr_pipe_0 <= addrb_2;
    end
    if (_GEN_96) begin
      mem_3__T_559_addr_pipe_0 <= addrb_3;
    end
    _T_74 <= rend;
    if (_T_74) begin
      _T_92_0 <= mem_0__T_61_data;
    end
    if (_T_74) begin
      _T_92_1 <= mem_1__T_61_data;
    end
    if (_T_74) begin
      _T_92_2 <= mem_2__T_61_data;
    end
    if (_T_74) begin
      _T_92_3 <= mem_3__T_61_data;
    end
    _T_329 <= renb;
    if (_T_329) begin
      _T_347_0 <= mem_0__T_316_data;
    end
    if (_T_329) begin
      _T_347_1 <= mem_1__T_316_data;
    end
    if (_T_329) begin
      _T_347_2 <= mem_2__T_316_data;
    end
    if (_T_329) begin
      _T_347_3 <= mem_3__T_316_data;
    end
    _T_410 <= renb;
    if (_T_410) begin
      _T_428_0 <= mem_0__T_397_data;
    end
    if (_T_410) begin
      _T_428_1 <= mem_1__T_397_data;
    end
    if (_T_410) begin
      _T_428_2 <= mem_2__T_397_data;
    end
    if (_T_410) begin
      _T_428_3 <= mem_3__T_397_data;
    end
    _T_491 <= renb;
    if (_T_491) begin
      _T_509_0 <= mem_0__T_478_data;
    end
    if (_T_491) begin
      _T_509_1 <= mem_1__T_478_data;
    end
    if (_T_491) begin
      _T_509_2 <= mem_2__T_478_data;
    end
    if (_T_491) begin
      _T_509_3 <= mem_3__T_478_data;
    end
    _T_572 <= renb;
    if (_T_572) begin
      _T_590_0 <= mem_0__T_559_data;
    end
    if (_T_572) begin
      _T_590_1 <= mem_1__T_559_data;
    end
    if (_T_572) begin
      _T_590_2 <= mem_2__T_559_data;
    end
    if (_T_572) begin
      _T_590_3 <= mem_3__T_559_data;
    end
  end
endmodule
module randomgen( // @[:@298.2]
  input         clock, // @[:@299.4]
  input         reset, // @[:@300.4]
  output [63:0] io_out, // @[:@301.4]
  input         io_en, // @[:@301.4]
  output        io_done // @[:@301.4]
);
  reg [63:0] curReg; // @[Random.scala 14:23:@303.4]
  reg [63:0] _RAND_0;
  reg [1:0] cnt; // @[Random.scala 15:20:@304.4]
  reg [31:0] _RAND_1;
  reg [15:0] _T_25; // @[LFSR.scala 22:23:@316.6]
  reg [31:0] _RAND_2;
  wire  _T_14; // @[Random.scala 19:28:@307.4]
  wire  _T_16; // @[Random.scala 19:17:@308.4]
  wire [2:0] _T_18; // @[Random.scala 22:23:@311.4]
  wire [1:0] _T_19; // @[Random.scala 22:23:@312.4]
  wire [1:0] _T_21; // @[Random.scala 22:13:@313.4]
  wire  _T_26; // @[LFSR.scala 23:40:@318.8]
  wire  _T_27; // @[LFSR.scala 23:48:@319.8]
  wire  _T_28; // @[LFSR.scala 23:43:@320.8]
  wire  _T_29; // @[LFSR.scala 23:56:@321.8]
  wire  _T_30; // @[LFSR.scala 23:51:@322.8]
  wire  _T_31; // @[LFSR.scala 23:64:@323.8]
  wire  _T_32; // @[LFSR.scala 23:59:@324.8]
  wire [14:0] _T_33; // @[LFSR.scala 23:73:@325.8]
  wire [15:0] _T_34; // @[Cat.scala 30:58:@326.8]
  wire [94:0] _GEN_2; // @[Random.scala 28:22:@329.6]
  wire [94:0] _T_36; // @[Random.scala 28:22:@329.6]
  wire [94:0] _GEN_3; // @[Random.scala 28:30:@330.6]
  wire [94:0] _T_37; // @[Random.scala 28:30:@330.6]
  wire [94:0] _GEN_1; // @[Random.scala 26:3:@315.4]
  assign _T_14 = cnt == 2'h0; // @[Random.scala 19:28:@307.4]
  assign _T_16 = io_en ? _T_14 : 1'h0; // @[Random.scala 19:17:@308.4]
  assign _T_18 = cnt + 2'h1; // @[Random.scala 22:23:@311.4]
  assign _T_19 = _T_18[1:0]; // @[Random.scala 22:23:@312.4]
  assign _T_21 = io_en ? _T_19 : 2'h0; // @[Random.scala 22:13:@313.4]
  assign _T_26 = _T_25[0]; // @[LFSR.scala 23:40:@318.8]
  assign _T_27 = _T_25[2]; // @[LFSR.scala 23:48:@319.8]
  assign _T_28 = _T_26 ^ _T_27; // @[LFSR.scala 23:43:@320.8]
  assign _T_29 = _T_25[3]; // @[LFSR.scala 23:56:@321.8]
  assign _T_30 = _T_28 ^ _T_29; // @[LFSR.scala 23:51:@322.8]
  assign _T_31 = _T_25[5]; // @[LFSR.scala 23:64:@323.8]
  assign _T_32 = _T_30 ^ _T_31; // @[LFSR.scala 23:59:@324.8]
  assign _T_33 = _T_25[15:1]; // @[LFSR.scala 23:73:@325.8]
  assign _T_34 = {_T_32,_T_33}; // @[Cat.scala 30:58:@326.8]
  assign _GEN_2 = {{31'd0}, curReg}; // @[Random.scala 28:22:@329.6]
  assign _T_36 = _GEN_2 << 5'h10; // @[Random.scala 28:22:@329.6]
  assign _GEN_3 = {{79'd0}, _T_25}; // @[Random.scala 28:30:@330.6]
  assign _T_37 = _T_36 | _GEN_3; // @[Random.scala 28:30:@330.6]
  assign _GEN_1 = io_en ? _T_37 : {{31'd0}, curReg}; // @[Random.scala 26:3:@315.4]
  assign io_out = curReg;
  assign io_done = _T_16;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{$random}};
  curReg = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  cnt = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  _T_25 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      curReg <= 64'h0;
    end else begin
      curReg <= _GEN_1[63:0];
    end
    if (reset) begin
      cnt <= 2'h0;
    end else begin
      if (io_en) begin
        cnt <= _T_19;
      end else begin
        cnt <= 2'h0;
      end
    end
    if (reset) begin
      _T_25 <= 16'h1;
    end else begin
      _T_25 <= _T_34;
    end
  end
endmodule
module counter( // @[:@334.2]
  input         clock, // @[:@335.4]
  input         io_get, // @[:@337.4]
  output [63:0] io_out, // @[:@337.4]
  input         io_reset, // @[:@337.4]
  input  [63:0] io_init // @[:@337.4]
);
  reg [63:0] cReg; // @[Counter.scala 15:17:@339.4]
  reg [63:0] _RAND_0;
  wire [64:0] _T_8; // @[Counter.scala 20:18:@340.4]
  wire [63:0] crp; // @[Counter.scala 20:18:@341.4]
  wire [63:0] _T_9; // @[Counter.scala 21:39:@342.4]
  wire [63:0] crp2; // @[Counter.scala 21:18:@343.4]
  wire  _T_10; // @[Counter.scala 28:15:@345.4]
  wire [63:0] _GEN_0; // @[Counter.scala 29:3:@346.4]
  assign _T_8 = cReg + 64'h1; // @[Counter.scala 20:18:@340.4]
  assign crp = _T_8[63:0]; // @[Counter.scala 20:18:@341.4]
  assign _T_9 = io_get ? crp : cReg; // @[Counter.scala 21:39:@342.4]
  assign crp2 = io_reset ? io_init : _T_9; // @[Counter.scala 21:18:@343.4]
  assign _T_10 = io_get | io_reset; // @[Counter.scala 28:15:@345.4]
  assign _GEN_0 = _T_10 ? crp2 : cReg; // @[Counter.scala 29:3:@346.4]
  assign io_out = crp2;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{$random}};
  cReg = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_10) begin
      if (io_reset) begin
        cReg <= io_init;
      end else begin
        if (io_get) begin
          cReg <= crp;
        end
      end
    end
  end
endmodule
module ivFileMac( // @[:@350.2]
  input          clock, // @[:@351.4]
  input          reset, // @[:@352.4]
  output [127:0] io_rdata, // @[:@353.4]
  input  [256:0] io_wdata, // @[:@353.4]
  input  [4:0]   io_addr, // @[:@353.4]
  input  [2:0]   io_cmd // @[:@353.4]
);
  reg [128:0] regmap_0; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_0;
  reg [128:0] regmap_1; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_1;
  reg [128:0] regmap_2; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_2;
  reg [128:0] regmap_3; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_3;
  reg [128:0] regmap_4; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_4;
  reg [128:0] regmap_5; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_5;
  reg [128:0] regmap_6; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_6;
  reg [128:0] regmap_7; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_7;
  reg [128:0] regmap_8; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_8;
  reg [128:0] regmap_9; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_9;
  reg [128:0] regmap_10; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_10;
  reg [128:0] regmap_11; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_11;
  reg [128:0] regmap_12; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_12;
  reg [128:0] regmap_13; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_13;
  reg [128:0] regmap_14; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_14;
  reg [128:0] regmap_15; // @[ivFileMac.scala 42:20:@372.4]
  reg [159:0] _RAND_15;
  reg [127:0] macreg_0; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_16;
  reg [127:0] macreg_1; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_17;
  reg [127:0] macreg_2; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_18;
  reg [127:0] macreg_3; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_19;
  reg [127:0] macreg_4; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_20;
  reg [127:0] macreg_5; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_21;
  reg [127:0] macreg_6; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_22;
  reg [127:0] macreg_7; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_23;
  reg [127:0] macreg_8; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_24;
  reg [127:0] macreg_9; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_25;
  reg [127:0] macreg_10; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_26;
  reg [127:0] macreg_11; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_27;
  reg [127:0] macreg_12; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_28;
  reg [127:0] macreg_13; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_29;
  reg [127:0] macreg_14; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_30;
  reg [127:0] macreg_15; // @[ivFileMac.scala 43:20:@390.4]
  reg [127:0] _RAND_31;
  reg [127:0] lastOut; // @[ivFileMac.scala 45:24:@391.4]
  reg [127:0] _RAND_32;
  wire  _T_260; // @[ivFileMac.scala 59:27:@394.4]
  wire  _T_262; // @[ivFileMac.scala 59:38:@395.4]
  wire  _T_264; // @[ivFileMac.scala 60:38:@396.4]
  wire  _T_266; // @[ivFileMac.scala 60:49:@397.4]
  wire  _T_268; // @[ivFileMac.scala 61:38:@398.4]
  wire  _T_270; // @[ivFileMac.scala 61:49:@399.4]
  wire  _T_272; // @[ivFileMac.scala 62:38:@400.4]
  wire  _T_274; // @[ivFileMac.scala 62:49:@401.4]
  wire  _T_276; // @[ivFileMac.scala 63:38:@402.4]
  wire  _T_278; // @[ivFileMac.scala 63:49:@403.4]
  wire  _T_280; // @[ivFileMac.scala 64:38:@404.4]
  wire  _T_282; // @[ivFileMac.scala 64:49:@405.4]
  wire  _T_284; // @[ivFileMac.scala 65:38:@406.4]
  wire  _T_286; // @[ivFileMac.scala 65:49:@407.4]
  wire  _T_288; // @[ivFileMac.scala 66:38:@408.4]
  wire  _T_290; // @[ivFileMac.scala 66:49:@409.4]
  wire  _T_292; // @[ivFileMac.scala 67:38:@410.4]
  wire  _T_294; // @[ivFileMac.scala 67:49:@411.4]
  wire  _T_296; // @[ivFileMac.scala 68:38:@412.4]
  wire  _T_298; // @[ivFileMac.scala 68:49:@413.4]
  wire  _T_300; // @[ivFileMac.scala 69:39:@414.4]
  wire  _T_302; // @[ivFileMac.scala 69:50:@415.4]
  wire  _T_304; // @[ivFileMac.scala 70:39:@416.4]
  wire  _T_306; // @[ivFileMac.scala 70:50:@417.4]
  wire  _T_308; // @[ivFileMac.scala 71:39:@418.4]
  wire  _T_310; // @[ivFileMac.scala 71:50:@419.4]
  wire  _T_312; // @[ivFileMac.scala 72:39:@420.4]
  wire  _T_314; // @[ivFileMac.scala 72:50:@421.4]
  wire  _T_316; // @[ivFileMac.scala 73:39:@422.4]
  wire  _T_318; // @[ivFileMac.scala 73:50:@423.4]
  wire  _T_320; // @[ivFileMac.scala 74:39:@424.4]
  wire  _T_322; // @[ivFileMac.scala 74:50:@425.4]
  wire [4:0] _T_325; // @[ivFileMac.scala 74:27:@426.4]
  wire [4:0] _T_326; // @[ivFileMac.scala 73:27:@427.4]
  wire [4:0] _T_327; // @[ivFileMac.scala 72:27:@428.4]
  wire [4:0] _T_328; // @[ivFileMac.scala 71:27:@429.4]
  wire [4:0] _T_329; // @[ivFileMac.scala 70:27:@430.4]
  wire [4:0] _T_330; // @[ivFileMac.scala 69:27:@431.4]
  wire [4:0] _T_331; // @[ivFileMac.scala 68:27:@432.4]
  wire [4:0] _T_332; // @[ivFileMac.scala 67:27:@433.4]
  wire [4:0] _T_333; // @[ivFileMac.scala 66:27:@434.4]
  wire [4:0] _T_334; // @[ivFileMac.scala 65:27:@435.4]
  wire [4:0] _T_335; // @[ivFileMac.scala 64:27:@436.4]
  wire [4:0] _T_336; // @[ivFileMac.scala 63:27:@437.4]
  wire [4:0] _T_337; // @[ivFileMac.scala 62:27:@438.4]
  wire [4:0] _T_338; // @[ivFileMac.scala 61:27:@439.4]
  wire [4:0] _T_339; // @[ivFileMac.scala 60:27:@440.4]
  wire [4:0] num; // @[ivFileMac.scala 59:16:@441.4]
  wire  _T_342; // @[ivFileMac.scala 83:30:@442.4]
  wire [3:0] _T_346; // @[:@443.4]
  wire [128:0] _GEN_6; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_7; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_8; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_9; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_10; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_11; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_12; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_13; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_14; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_15; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_16; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_17; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_18; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_19; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _GEN_20; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_21; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_22; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_23; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_24; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_25; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_26; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_27; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_28; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_29; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_30; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_31; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_32; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_33; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_34; // @[ivFileMac.scala 83:21:@445.4]
  wire [127:0] _GEN_35; // @[ivFileMac.scala 83:21:@445.4]
  wire [128:0] _T_351; // @[ivFileMac.scala 83:21:@445.4]
  wire  _T_358; // @[Mux.scala 46:19:@447.4]
  wire [127:0] _T_359; // @[Mux.scala 46:16:@448.4]
  wire  _T_360; // @[Mux.scala 46:19:@449.4]
  wire [127:0] _T_361; // @[Mux.scala 46:16:@450.4]
  wire  _T_362; // @[Mux.scala 46:19:@451.4]
  wire [128:0] rout; // @[Mux.scala 46:16:@452.4]
  wire  _T_364; // @[ivFileMac.scala 88:24:@453.4]
  wire  _T_366; // @[ivFileMac.scala 88:42:@454.4]
  wire  _T_367; // @[ivFileMac.scala 88:32:@455.4]
  wire  _T_369; // @[ivFileMac.scala 88:60:@456.4]
  wire  cmdRead; // @[ivFileMac.scala 88:50:@457.4]
  wire [128:0] _T_370; // @[ivFileMac.scala 91:17:@459.4]
  wire  _T_372; // @[ivFileMac.scala 100:17:@461.4]
  wire [128:0] _T_373; // @[ivFileMac.scala 102:33:@463.6]
  wire [127:0] _T_374; // @[ivFileMac.scala 103:32:@464.6]
  wire [128:0] _GEN_51; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_52; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_53; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_54; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_55; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_56; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_57; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_58; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_59; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_60; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_61; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_62; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_63; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_64; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_65; // @[ivFileMac.scala 107:27:@468.8]
  wire [128:0] _GEN_66; // @[ivFileMac.scala 107:27:@468.8]
  wire [127:0] _GEN_67; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_68; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_69; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_70; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_71; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_72; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_73; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_74; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_75; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_76; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_77; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_78; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_79; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_80; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_81; // @[ivFileMac.scala 108:27:@470.8]
  wire [127:0] _GEN_82; // @[ivFileMac.scala 108:27:@470.8]
  wire [128:0] _GEN_99; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_100; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_101; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_102; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_103; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_104; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_105; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_106; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_107; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_108; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_109; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_110; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_111; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_112; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_113; // @[ivFileMac.scala 106:9:@466.6]
  wire [128:0] _GEN_114; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_115; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_116; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_117; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_118; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_119; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_120; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_121; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_122; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_123; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_124; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_125; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_126; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_127; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_128; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_129; // @[ivFileMac.scala 106:9:@466.6]
  wire [127:0] _GEN_130; // @[ivFileMac.scala 106:9:@466.6]
  wire  _T_390; // @[ivFileMac.scala 115:23:@478.6]
  wire [112:0] _GEN_131; // @[ivFileMac.scala 116:5:@479.6]
  wire [125:0] _GEN_132; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_133; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_134; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_135; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_136; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_137; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_138; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_139; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_140; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_141; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_142; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_143; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_144; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_145; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_146; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_147; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_148; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_149; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_150; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_151; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_152; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_153; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_154; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_155; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_156; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_157; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_158; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_159; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_160; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_161; // @[ivFileMac.scala 116:5:@479.6]
  wire [127:0] _GEN_162; // @[ivFileMac.scala 116:5:@479.6]
  wire [128:0] _GEN_163; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_164; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_165; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_166; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_167; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_168; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_169; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_170; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_171; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_172; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_173; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_174; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_175; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_176; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_177; // @[ivFileMac.scala 101:5:@462.4]
  wire [128:0] _GEN_178; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_179; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_180; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_181; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_182; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_183; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_184; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_185; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_186; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_187; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_188; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_189; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_190; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_191; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_192; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_193; // @[ivFileMac.scala 101:5:@462.4]
  wire [127:0] _GEN_194; // @[ivFileMac.scala 101:5:@462.4]
  assign _T_260 = regmap_0[128]; // @[ivFileMac.scala 59:27:@394.4]
  assign _T_262 = _T_260 == 1'h0; // @[ivFileMac.scala 59:38:@395.4]
  assign _T_264 = regmap_1[128]; // @[ivFileMac.scala 60:38:@396.4]
  assign _T_266 = _T_264 == 1'h0; // @[ivFileMac.scala 60:49:@397.4]
  assign _T_268 = regmap_2[128]; // @[ivFileMac.scala 61:38:@398.4]
  assign _T_270 = _T_268 == 1'h0; // @[ivFileMac.scala 61:49:@399.4]
  assign _T_272 = regmap_3[128]; // @[ivFileMac.scala 62:38:@400.4]
  assign _T_274 = _T_272 == 1'h0; // @[ivFileMac.scala 62:49:@401.4]
  assign _T_276 = regmap_4[128]; // @[ivFileMac.scala 63:38:@402.4]
  assign _T_278 = _T_276 == 1'h0; // @[ivFileMac.scala 63:49:@403.4]
  assign _T_280 = regmap_5[128]; // @[ivFileMac.scala 64:38:@404.4]
  assign _T_282 = _T_280 == 1'h0; // @[ivFileMac.scala 64:49:@405.4]
  assign _T_284 = regmap_6[128]; // @[ivFileMac.scala 65:38:@406.4]
  assign _T_286 = _T_284 == 1'h0; // @[ivFileMac.scala 65:49:@407.4]
  assign _T_288 = regmap_7[128]; // @[ivFileMac.scala 66:38:@408.4]
  assign _T_290 = _T_288 == 1'h0; // @[ivFileMac.scala 66:49:@409.4]
  assign _T_292 = regmap_8[128]; // @[ivFileMac.scala 67:38:@410.4]
  assign _T_294 = _T_292 == 1'h0; // @[ivFileMac.scala 67:49:@411.4]
  assign _T_296 = regmap_9[128]; // @[ivFileMac.scala 68:38:@412.4]
  assign _T_298 = _T_296 == 1'h0; // @[ivFileMac.scala 68:49:@413.4]
  assign _T_300 = regmap_10[128]; // @[ivFileMac.scala 69:39:@414.4]
  assign _T_302 = _T_300 == 1'h0; // @[ivFileMac.scala 69:50:@415.4]
  assign _T_304 = regmap_11[128]; // @[ivFileMac.scala 70:39:@416.4]
  assign _T_306 = _T_304 == 1'h0; // @[ivFileMac.scala 70:50:@417.4]
  assign _T_308 = regmap_12[128]; // @[ivFileMac.scala 71:39:@418.4]
  assign _T_310 = _T_308 == 1'h0; // @[ivFileMac.scala 71:50:@419.4]
  assign _T_312 = regmap_13[128]; // @[ivFileMac.scala 72:39:@420.4]
  assign _T_314 = _T_312 == 1'h0; // @[ivFileMac.scala 72:50:@421.4]
  assign _T_316 = regmap_14[128]; // @[ivFileMac.scala 73:39:@422.4]
  assign _T_318 = _T_316 == 1'h0; // @[ivFileMac.scala 73:50:@423.4]
  assign _T_320 = regmap_15[128]; // @[ivFileMac.scala 74:39:@424.4]
  assign _T_322 = _T_320 == 1'h0; // @[ivFileMac.scala 74:50:@425.4]
  assign _T_325 = _T_322 ? 5'hf : 5'h10; // @[ivFileMac.scala 74:27:@426.4]
  assign _T_326 = _T_318 ? 5'he : _T_325; // @[ivFileMac.scala 73:27:@427.4]
  assign _T_327 = _T_314 ? 5'hd : _T_326; // @[ivFileMac.scala 72:27:@428.4]
  assign _T_328 = _T_310 ? 5'hc : _T_327; // @[ivFileMac.scala 71:27:@429.4]
  assign _T_329 = _T_306 ? 5'hb : _T_328; // @[ivFileMac.scala 70:27:@430.4]
  assign _T_330 = _T_302 ? 5'ha : _T_329; // @[ivFileMac.scala 69:27:@431.4]
  assign _T_331 = _T_298 ? 5'h9 : _T_330; // @[ivFileMac.scala 68:27:@432.4]
  assign _T_332 = _T_294 ? 5'h8 : _T_331; // @[ivFileMac.scala 67:27:@433.4]
  assign _T_333 = _T_290 ? 5'h7 : _T_332; // @[ivFileMac.scala 66:27:@434.4]
  assign _T_334 = _T_286 ? 5'h6 : _T_333; // @[ivFileMac.scala 65:27:@435.4]
  assign _T_335 = _T_282 ? 5'h5 : _T_334; // @[ivFileMac.scala 64:27:@436.4]
  assign _T_336 = _T_278 ? 5'h4 : _T_335; // @[ivFileMac.scala 63:27:@437.4]
  assign _T_337 = _T_274 ? 5'h3 : _T_336; // @[ivFileMac.scala 62:27:@438.4]
  assign _T_338 = _T_270 ? 5'h2 : _T_337; // @[ivFileMac.scala 61:27:@439.4]
  assign _T_339 = _T_266 ? 5'h1 : _T_338; // @[ivFileMac.scala 60:27:@440.4]
  assign num = _T_262 ? 5'h0 : _T_339; // @[ivFileMac.scala 59:16:@441.4]
  assign _T_342 = io_addr <= 5'hf; // @[ivFileMac.scala 83:30:@442.4]
  assign _T_346 = io_addr[3:0]; // @[:@443.4]
  assign _GEN_6 = 4'h1 == _T_346 ? regmap_1 : regmap_0; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_7 = 4'h2 == _T_346 ? regmap_2 : _GEN_6; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_8 = 4'h3 == _T_346 ? regmap_3 : _GEN_7; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_9 = 4'h4 == _T_346 ? regmap_4 : _GEN_8; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_10 = 4'h5 == _T_346 ? regmap_5 : _GEN_9; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_11 = 4'h6 == _T_346 ? regmap_6 : _GEN_10; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_12 = 4'h7 == _T_346 ? regmap_7 : _GEN_11; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_13 = 4'h8 == _T_346 ? regmap_8 : _GEN_12; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_14 = 4'h9 == _T_346 ? regmap_9 : _GEN_13; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_15 = 4'ha == _T_346 ? regmap_10 : _GEN_14; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_16 = 4'hb == _T_346 ? regmap_11 : _GEN_15; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_17 = 4'hc == _T_346 ? regmap_12 : _GEN_16; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_18 = 4'hd == _T_346 ? regmap_13 : _GEN_17; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_19 = 4'he == _T_346 ? regmap_14 : _GEN_18; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_20 = 4'hf == _T_346 ? regmap_15 : _GEN_19; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_21 = 4'h1 == _T_346 ? macreg_1 : macreg_0; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_22 = 4'h2 == _T_346 ? macreg_2 : _GEN_21; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_23 = 4'h3 == _T_346 ? macreg_3 : _GEN_22; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_24 = 4'h4 == _T_346 ? macreg_4 : _GEN_23; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_25 = 4'h5 == _T_346 ? macreg_5 : _GEN_24; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_26 = 4'h6 == _T_346 ? macreg_6 : _GEN_25; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_27 = 4'h7 == _T_346 ? macreg_7 : _GEN_26; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_28 = 4'h8 == _T_346 ? macreg_8 : _GEN_27; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_29 = 4'h9 == _T_346 ? macreg_9 : _GEN_28; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_30 = 4'ha == _T_346 ? macreg_10 : _GEN_29; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_31 = 4'hb == _T_346 ? macreg_11 : _GEN_30; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_32 = 4'hc == _T_346 ? macreg_12 : _GEN_31; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_33 = 4'hd == _T_346 ? macreg_13 : _GEN_32; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_34 = 4'he == _T_346 ? macreg_14 : _GEN_33; // @[ivFileMac.scala 83:21:@445.4]
  assign _GEN_35 = 4'hf == _T_346 ? macreg_15 : _GEN_34; // @[ivFileMac.scala 83:21:@445.4]
  assign _T_351 = _T_342 ? _GEN_20 : {{1'd0}, _GEN_35}; // @[ivFileMac.scala 83:21:@445.4]
  assign _T_358 = 3'h6 == io_cmd; // @[Mux.scala 46:19:@447.4]
  assign _T_359 = _T_358 ? {{123'd0}, num} : lastOut; // @[Mux.scala 46:16:@448.4]
  assign _T_360 = 3'h3 == io_cmd; // @[Mux.scala 46:19:@449.4]
  assign _T_361 = _T_360 ? _GEN_35 : _T_359; // @[Mux.scala 46:16:@450.4]
  assign _T_362 = 3'h1 == io_cmd; // @[Mux.scala 46:19:@451.4]
  assign rout = _T_362 ? _T_351 : {{1'd0}, _T_361}; // @[Mux.scala 46:16:@452.4]
  assign _T_364 = io_cmd == 3'h1; // @[ivFileMac.scala 88:24:@453.4]
  assign _T_366 = io_cmd == 3'h3; // @[ivFileMac.scala 88:42:@454.4]
  assign _T_367 = _T_364 | _T_366; // @[ivFileMac.scala 88:32:@455.4]
  assign _T_369 = io_cmd == 3'h6; // @[ivFileMac.scala 88:60:@456.4]
  assign cmdRead = _T_367 | _T_369; // @[ivFileMac.scala 88:50:@457.4]
  assign _T_370 = cmdRead ? rout : {{1'd0}, lastOut}; // @[ivFileMac.scala 91:17:@459.4]
  assign _T_372 = io_cmd == 3'h2; // @[ivFileMac.scala 100:17:@461.4]
  assign _T_373 = io_wdata[256:128]; // @[ivFileMac.scala 102:33:@463.6]
  assign _T_374 = io_wdata[127:0]; // @[ivFileMac.scala 103:32:@464.6]
  assign _GEN_51 = 4'h0 == _T_346 ? _T_373 : 129'h180004000200080104008a004d002; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_52 = 4'h1 == _T_346 ? _T_373 : regmap_1; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_53 = 4'h2 == _T_346 ? _T_373 : regmap_2; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_54 = 4'h3 == _T_346 ? _T_373 : regmap_3; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_55 = 4'h4 == _T_346 ? _T_373 : regmap_4; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_56 = 4'h5 == _T_346 ? _T_373 : regmap_5; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_57 = 4'h6 == _T_346 ? _T_373 : regmap_6; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_58 = 4'h7 == _T_346 ? _T_373 : regmap_7; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_59 = 4'h8 == _T_346 ? _T_373 : regmap_8; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_60 = 4'h9 == _T_346 ? _T_373 : regmap_9; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_61 = 4'ha == _T_346 ? _T_373 : regmap_10; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_62 = 4'hb == _T_346 ? _T_373 : regmap_11; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_63 = 4'hc == _T_346 ? _T_373 : regmap_12; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_64 = 4'hd == _T_346 ? _T_373 : regmap_13; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_65 = 4'he == _T_346 ? _T_373 : regmap_14; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_66 = 4'hf == _T_346 ? _T_373 : regmap_15; // @[ivFileMac.scala 107:27:@468.8]
  assign _GEN_67 = 4'h0 == _T_346 ? _T_374 : 128'h3de39d24188a846a636f37b0f69124e6; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_68 = 4'h1 == _T_346 ? _T_374 : macreg_1; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_69 = 4'h2 == _T_346 ? _T_374 : macreg_2; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_70 = 4'h3 == _T_346 ? _T_374 : macreg_3; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_71 = 4'h4 == _T_346 ? _T_374 : macreg_4; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_72 = 4'h5 == _T_346 ? _T_374 : macreg_5; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_73 = 4'h6 == _T_346 ? _T_374 : macreg_6; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_74 = 4'h7 == _T_346 ? _T_374 : macreg_7; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_75 = 4'h8 == _T_346 ? _T_374 : macreg_8; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_76 = 4'h9 == _T_346 ? _T_374 : macreg_9; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_77 = 4'ha == _T_346 ? _T_374 : macreg_10; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_78 = 4'hb == _T_346 ? _T_374 : macreg_11; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_79 = 4'hc == _T_346 ? _T_374 : macreg_12; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_80 = 4'hd == _T_346 ? _T_374 : macreg_13; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_81 = 4'he == _T_346 ? _T_374 : macreg_14; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_82 = 4'hf == _T_346 ? _T_374 : macreg_15; // @[ivFileMac.scala 108:27:@470.8]
  assign _GEN_99 = _T_342 ? _GEN_51 : 129'h180004000200080104008a004d002; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_100 = _T_342 ? _GEN_52 : regmap_1; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_101 = _T_342 ? _GEN_53 : regmap_2; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_102 = _T_342 ? _GEN_54 : regmap_3; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_103 = _T_342 ? _GEN_55 : regmap_4; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_104 = _T_342 ? _GEN_56 : regmap_5; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_105 = _T_342 ? _GEN_57 : regmap_6; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_106 = _T_342 ? _GEN_58 : regmap_7; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_107 = _T_342 ? _GEN_59 : regmap_8; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_108 = _T_342 ? _GEN_60 : regmap_9; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_109 = _T_342 ? _GEN_61 : regmap_10; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_110 = _T_342 ? _GEN_62 : regmap_11; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_111 = _T_342 ? _GEN_63 : regmap_12; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_112 = _T_342 ? _GEN_64 : regmap_13; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_113 = _T_342 ? _GEN_65 : regmap_14; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_114 = _T_342 ? _GEN_66 : regmap_15; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_115 = _T_342 ? _GEN_67 : _GEN_67; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_116 = _T_342 ? _GEN_68 : _GEN_68; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_117 = _T_342 ? _GEN_69 : _GEN_69; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_118 = _T_342 ? _GEN_70 : _GEN_70; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_119 = _T_342 ? _GEN_71 : _GEN_71; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_120 = _T_342 ? _GEN_72 : _GEN_72; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_121 = _T_342 ? _GEN_73 : _GEN_73; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_122 = _T_342 ? _GEN_74 : _GEN_74; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_123 = _T_342 ? _GEN_75 : _GEN_75; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_124 = _T_342 ? _GEN_76 : _GEN_76; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_125 = _T_342 ? _GEN_77 : _GEN_77; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_126 = _T_342 ? _GEN_78 : _GEN_78; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_127 = _T_342 ? _GEN_79 : _GEN_79; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_128 = _T_342 ? _GEN_80 : _GEN_80; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_129 = _T_342 ? _GEN_81 : _GEN_81; // @[ivFileMac.scala 106:9:@466.6]
  assign _GEN_130 = _T_342 ? _GEN_82 : _GEN_82; // @[ivFileMac.scala 106:9:@466.6]
  assign _T_390 = io_cmd == 3'h5; // @[ivFileMac.scala 115:23:@478.6]
  assign _GEN_131 = _T_390 ? 113'h0 : 113'h180004000200080104008a004d002; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_132 = _T_390 ? 126'h0 : 126'h3de39d24188a846a636f37b0f69124e6; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_133 = _T_390 ? 129'h0 : regmap_1; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_134 = _T_390 ? 128'h0 : macreg_1; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_135 = _T_390 ? 129'h0 : regmap_2; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_136 = _T_390 ? 128'h0 : macreg_2; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_137 = _T_390 ? 129'h0 : regmap_3; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_138 = _T_390 ? 128'h0 : macreg_3; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_139 = _T_390 ? 129'h0 : regmap_4; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_140 = _T_390 ? 128'h0 : macreg_4; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_141 = _T_390 ? 129'h0 : regmap_5; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_142 = _T_390 ? 128'h0 : macreg_5; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_143 = _T_390 ? 129'h0 : regmap_6; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_144 = _T_390 ? 128'h0 : macreg_6; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_145 = _T_390 ? 129'h0 : regmap_7; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_146 = _T_390 ? 128'h0 : macreg_7; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_147 = _T_390 ? 129'h0 : regmap_8; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_148 = _T_390 ? 128'h0 : macreg_8; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_149 = _T_390 ? 129'h0 : regmap_9; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_150 = _T_390 ? 128'h0 : macreg_9; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_151 = _T_390 ? 129'h0 : regmap_10; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_152 = _T_390 ? 128'h0 : macreg_10; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_153 = _T_390 ? 129'h0 : regmap_11; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_154 = _T_390 ? 128'h0 : macreg_11; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_155 = _T_390 ? 129'h0 : regmap_12; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_156 = _T_390 ? 128'h0 : macreg_12; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_157 = _T_390 ? 129'h0 : regmap_13; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_158 = _T_390 ? 128'h0 : macreg_13; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_159 = _T_390 ? 129'h0 : regmap_14; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_160 = _T_390 ? 128'h0 : macreg_14; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_161 = _T_390 ? 129'h0 : regmap_15; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_162 = _T_390 ? 128'h0 : macreg_15; // @[ivFileMac.scala 116:5:@479.6]
  assign _GEN_163 = _T_372 ? _GEN_99 : {{16'd0}, _GEN_131}; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_164 = _T_372 ? _GEN_100 : _GEN_133; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_165 = _T_372 ? _GEN_101 : _GEN_135; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_166 = _T_372 ? _GEN_102 : _GEN_137; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_167 = _T_372 ? _GEN_103 : _GEN_139; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_168 = _T_372 ? _GEN_104 : _GEN_141; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_169 = _T_372 ? _GEN_105 : _GEN_143; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_170 = _T_372 ? _GEN_106 : _GEN_145; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_171 = _T_372 ? _GEN_107 : _GEN_147; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_172 = _T_372 ? _GEN_108 : _GEN_149; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_173 = _T_372 ? _GEN_109 : _GEN_151; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_174 = _T_372 ? _GEN_110 : _GEN_153; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_175 = _T_372 ? _GEN_111 : _GEN_155; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_176 = _T_372 ? _GEN_112 : _GEN_157; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_177 = _T_372 ? _GEN_113 : _GEN_159; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_178 = _T_372 ? _GEN_114 : _GEN_161; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_179 = _T_372 ? _GEN_115 : {{2'd0}, _GEN_132}; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_180 = _T_372 ? _GEN_116 : _GEN_134; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_181 = _T_372 ? _GEN_117 : _GEN_136; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_182 = _T_372 ? _GEN_118 : _GEN_138; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_183 = _T_372 ? _GEN_119 : _GEN_140; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_184 = _T_372 ? _GEN_120 : _GEN_142; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_185 = _T_372 ? _GEN_121 : _GEN_144; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_186 = _T_372 ? _GEN_122 : _GEN_146; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_187 = _T_372 ? _GEN_123 : _GEN_148; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_188 = _T_372 ? _GEN_124 : _GEN_150; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_189 = _T_372 ? _GEN_125 : _GEN_152; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_190 = _T_372 ? _GEN_126 : _GEN_154; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_191 = _T_372 ? _GEN_127 : _GEN_156; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_192 = _T_372 ? _GEN_128 : _GEN_158; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_193 = _T_372 ? _GEN_129 : _GEN_160; // @[ivFileMac.scala 101:5:@462.4]
  assign _GEN_194 = _T_372 ? _GEN_130 : _GEN_162; // @[ivFileMac.scala 101:5:@462.4]
  assign io_rdata = rout[127:0];
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{$random}};
  regmap_0 = _RAND_0[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {5{$random}};
  regmap_1 = _RAND_1[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {5{$random}};
  regmap_2 = _RAND_2[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {5{$random}};
  regmap_3 = _RAND_3[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {5{$random}};
  regmap_4 = _RAND_4[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {5{$random}};
  regmap_5 = _RAND_5[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {5{$random}};
  regmap_6 = _RAND_6[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {5{$random}};
  regmap_7 = _RAND_7[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {5{$random}};
  regmap_8 = _RAND_8[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {5{$random}};
  regmap_9 = _RAND_9[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {5{$random}};
  regmap_10 = _RAND_10[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {5{$random}};
  regmap_11 = _RAND_11[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {5{$random}};
  regmap_12 = _RAND_12[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {5{$random}};
  regmap_13 = _RAND_13[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {5{$random}};
  regmap_14 = _RAND_14[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {5{$random}};
  regmap_15 = _RAND_15[128:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {4{$random}};
  macreg_0 = _RAND_16[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {4{$random}};
  macreg_1 = _RAND_17[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {4{$random}};
  macreg_2 = _RAND_18[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {4{$random}};
  macreg_3 = _RAND_19[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {4{$random}};
  macreg_4 = _RAND_20[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {4{$random}};
  macreg_5 = _RAND_21[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {4{$random}};
  macreg_6 = _RAND_22[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {4{$random}};
  macreg_7 = _RAND_23[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {4{$random}};
  macreg_8 = _RAND_24[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {4{$random}};
  macreg_9 = _RAND_25[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {4{$random}};
  macreg_10 = _RAND_26[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {4{$random}};
  macreg_11 = _RAND_27[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {4{$random}};
  macreg_12 = _RAND_28[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {4{$random}};
  macreg_13 = _RAND_29[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {4{$random}};
  macreg_14 = _RAND_30[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {4{$random}};
  macreg_15 = _RAND_31[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {4{$random}};
  lastOut = _RAND_32[127:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regmap_0 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h0 == _T_346) begin
            regmap_0 <= _T_373;
          end else begin
            regmap_0 <= 129'h180004000200080104008a004d002;
          end
        end else begin
          regmap_0 <= 129'h180004000200080104008a004d002;
        end
      end else begin
        regmap_0 <= {{16'd0}, _GEN_131};
      end
    end
    if (reset) begin
      regmap_1 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h1 == _T_346) begin
            regmap_1 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_1 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_2 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h2 == _T_346) begin
            regmap_2 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_2 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_3 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h3 == _T_346) begin
            regmap_3 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_3 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_4 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h4 == _T_346) begin
            regmap_4 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_4 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_5 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h5 == _T_346) begin
            regmap_5 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_5 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_6 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h6 == _T_346) begin
            regmap_6 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_6 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_7 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h7 == _T_346) begin
            regmap_7 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_7 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_8 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h8 == _T_346) begin
            regmap_8 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_8 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_9 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h9 == _T_346) begin
            regmap_9 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_9 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_10 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'ha == _T_346) begin
            regmap_10 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_10 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_11 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hb == _T_346) begin
            regmap_11 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_11 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_12 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hc == _T_346) begin
            regmap_12 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_12 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_13 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hd == _T_346) begin
            regmap_13 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_13 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_14 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'he == _T_346) begin
            regmap_14 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_14 <= 129'h0;
        end
      end
    end
    if (reset) begin
      regmap_15 <= 129'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hf == _T_346) begin
            regmap_15 <= _T_373;
          end
        end
      end else begin
        if (_T_390) begin
          regmap_15 <= 129'h0;
        end
      end
    end
    if (reset) begin
      macreg_0 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h0 == _T_346) begin
            macreg_0 <= _T_374;
          end else begin
            macreg_0 <= 128'h3de39d24188a846a636f37b0f69124e6;
          end
        end else begin
          if (4'h0 == _T_346) begin
            macreg_0 <= _T_374;
          end else begin
            macreg_0 <= 128'h3de39d24188a846a636f37b0f69124e6;
          end
        end
      end else begin
        macreg_0 <= {{2'd0}, _GEN_132};
      end
    end
    if (reset) begin
      macreg_1 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h1 == _T_346) begin
            macreg_1 <= _T_374;
          end
        end else begin
          if (4'h1 == _T_346) begin
            macreg_1 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_1 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_2 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h2 == _T_346) begin
            macreg_2 <= _T_374;
          end
        end else begin
          if (4'h2 == _T_346) begin
            macreg_2 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_2 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_3 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h3 == _T_346) begin
            macreg_3 <= _T_374;
          end
        end else begin
          if (4'h3 == _T_346) begin
            macreg_3 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_3 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_4 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h4 == _T_346) begin
            macreg_4 <= _T_374;
          end
        end else begin
          if (4'h4 == _T_346) begin
            macreg_4 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_4 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_5 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h5 == _T_346) begin
            macreg_5 <= _T_374;
          end
        end else begin
          if (4'h5 == _T_346) begin
            macreg_5 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_5 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_6 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h6 == _T_346) begin
            macreg_6 <= _T_374;
          end
        end else begin
          if (4'h6 == _T_346) begin
            macreg_6 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_6 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_7 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h7 == _T_346) begin
            macreg_7 <= _T_374;
          end
        end else begin
          if (4'h7 == _T_346) begin
            macreg_7 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_7 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_8 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h8 == _T_346) begin
            macreg_8 <= _T_374;
          end
        end else begin
          if (4'h8 == _T_346) begin
            macreg_8 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_8 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_9 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'h9 == _T_346) begin
            macreg_9 <= _T_374;
          end
        end else begin
          if (4'h9 == _T_346) begin
            macreg_9 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_9 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_10 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'ha == _T_346) begin
            macreg_10 <= _T_374;
          end
        end else begin
          if (4'ha == _T_346) begin
            macreg_10 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_10 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_11 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hb == _T_346) begin
            macreg_11 <= _T_374;
          end
        end else begin
          if (4'hb == _T_346) begin
            macreg_11 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_11 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_12 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hc == _T_346) begin
            macreg_12 <= _T_374;
          end
        end else begin
          if (4'hc == _T_346) begin
            macreg_12 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_12 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_13 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hd == _T_346) begin
            macreg_13 <= _T_374;
          end
        end else begin
          if (4'hd == _T_346) begin
            macreg_13 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_13 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_14 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'he == _T_346) begin
            macreg_14 <= _T_374;
          end
        end else begin
          if (4'he == _T_346) begin
            macreg_14 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_14 <= 128'h0;
        end
      end
    end
    if (reset) begin
      macreg_15 <= 128'h0;
    end else begin
      if (_T_372) begin
        if (_T_342) begin
          if (4'hf == _T_346) begin
            macreg_15 <= _T_374;
          end
        end else begin
          if (4'hf == _T_346) begin
            macreg_15 <= _T_374;
          end
        end
      end else begin
        if (_T_390) begin
          macreg_15 <= 128'h0;
        end
      end
    end
    if (reset) begin
      lastOut <= 128'h0;
    end else begin
      lastOut <= _T_370[127:0];
    end
  end
endmodule
module enc( // @[:@514.2]
  input          clock, // @[:@515.4]
  input          reset, // @[:@516.4]
  input  [127:0] io_rkey, // @[:@517.4]
  output         io_done, // @[:@517.4]
  output [127:0] io_sio_addr2, // @[:@517.4]
  input  [127:0] io_sio_data2, // @[:@517.4]
  output [127:0] io_out, // @[:@517.4]
  output [3:0]   io_roundOut, // @[:@517.4]
  input  [127:0] io_data, // @[:@517.4]
  input          io_en // @[:@517.4]
);
  reg [3:0] roundCounter; // @[aesencrypt.scala 22:29:@519.4]
  reg [31:0] _RAND_0;
  reg [127:0] state; // @[aesencrypt.scala 23:22:@520.4]
  reg [127:0] _RAND_1;
  wire  _T_19; // @[aesencrypt.scala 24:37:@521.4]
  wire  _T_21; // @[aesencrypt.scala 24:17:@522.4]
  wire [4:0] _T_23; // @[aesencrypt.scala 43:42:@524.4]
  wire [3:0] _T_24; // @[aesencrypt.scala 43:42:@525.4]
  wire [3:0] _T_26; // @[aesencrypt.scala 43:22:@526.4]
  wire [3:0] _T_28; // @[aesencrypt.scala 44:21:@528.4]
  wire [127:0] t; // @[aesencrypt.scala 156:25:@530.4]
  wire [7:0] _T_29; // @[aesencrypt.scala 168:14:@532.4]
  wire [7:0] _T_30; // @[aesencrypt.scala 169:14:@533.4]
  wire [7:0] _T_31; // @[aesencrypt.scala 170:14:@534.4]
  wire [7:0] _T_32; // @[aesencrypt.scala 171:14:@535.4]
  wire [15:0] _T_33; // @[Cat.scala 30:58:@536.4]
  wire [15:0] _T_34; // @[Cat.scala 30:58:@537.4]
  wire [31:0] _T_35; // @[Cat.scala 30:58:@538.4]
  wire [7:0] _T_36; // @[aesencrypt.scala 174:15:@539.4]
  wire [7:0] _T_37; // @[aesencrypt.scala 175:15:@540.4]
  wire [7:0] _T_38; // @[aesencrypt.scala 177:14:@541.4]
  wire [7:0] _T_39; // @[aesencrypt.scala 178:14:@542.4]
  wire [15:0] _T_40; // @[Cat.scala 30:58:@543.4]
  wire [15:0] _T_41; // @[Cat.scala 30:58:@544.4]
  wire [31:0] _T_42; // @[Cat.scala 30:58:@545.4]
  wire [7:0] _T_43; // @[aesencrypt.scala 181:15:@546.4]
  wire [7:0] _T_44; // @[aesencrypt.scala 182:15:@547.4]
  wire [7:0] _T_45; // @[aesencrypt.scala 183:15:@548.4]
  wire [7:0] _T_46; // @[aesencrypt.scala 184:15:@549.4]
  wire [15:0] _T_47; // @[Cat.scala 30:58:@550.4]
  wire [15:0] _T_48; // @[Cat.scala 30:58:@551.4]
  wire [31:0] _T_49; // @[Cat.scala 30:58:@552.4]
  wire [7:0] _T_50; // @[aesencrypt.scala 187:14:@553.4]
  wire [7:0] _T_51; // @[aesencrypt.scala 188:14:@554.4]
  wire [7:0] _T_52; // @[aesencrypt.scala 189:14:@555.4]
  wire [7:0] _T_53; // @[aesencrypt.scala 190:14:@556.4]
  wire [15:0] _T_54; // @[Cat.scala 30:58:@557.4]
  wire [15:0] _T_55; // @[Cat.scala 30:58:@558.4]
  wire [31:0] _T_56; // @[Cat.scala 30:58:@559.4]
  wire [63:0] _T_57; // @[Cat.scala 30:58:@560.4]
  wire [63:0] _T_58; // @[Cat.scala 30:58:@561.4]
  wire [127:0] state1; // @[Cat.scala 30:58:@562.4]
  wire [7:0] _T_59; // @[aesencrypt.scala 220:21:@563.4]
  wire [7:0] _T_60; // @[aesencrypt.scala 221:21:@564.4]
  wire [7:0] _T_61; // @[aesencrypt.scala 222:21:@565.4]
  wire [7:0] _T_62; // @[aesencrypt.scala 223:21:@566.4]
  wire [7:0] _T_63; // @[aesencrypt.scala 231:23:@567.4]
  wire [7:0] _T_64; // @[aesencrypt.scala 231:32:@568.4]
  wire [7:0] _T_65; // @[aesencrypt.scala 231:41:@569.4]
  wire [8:0] _GEN_10; // @[aesencrypt.scala 198:27:@571.4]
  wire [8:0] _T_68; // @[aesencrypt.scala 198:27:@571.4]
  wire [8:0] _T_70; // @[aesencrypt.scala 198:35:@572.4]
  wire [7:0] _T_71; // @[aesencrypt.scala 198:46:@573.4]
  wire [7:0] _T_74; // @[aesencrypt.scala 199:31:@575.4]
  wire [7:0] _T_76; // @[aesencrypt.scala 200:25:@576.4]
  wire  _T_78; // @[aesencrypt.scala 200:36:@577.4]
  wire [7:0] _T_79; // @[aesencrypt.scala 201:18:@578.4]
  wire [7:0] _T_80; // @[aesencrypt.scala 238:25:@579.4]
  wire [7:0] _T_81; // @[aesencrypt.scala 238:32:@580.4]
  wire [7:0] _T_82; // @[aesencrypt.scala 241:26:@581.4]
  wire [8:0] _GEN_12; // @[aesencrypt.scala 198:27:@582.4]
  wire [8:0] _T_84; // @[aesencrypt.scala 198:27:@582.4]
  wire [8:0] _T_86; // @[aesencrypt.scala 198:35:@583.4]
  wire [7:0] _T_87; // @[aesencrypt.scala 198:46:@584.4]
  wire [7:0] _T_90; // @[aesencrypt.scala 199:31:@586.4]
  wire [7:0] _T_92; // @[aesencrypt.scala 200:25:@587.4]
  wire  _T_94; // @[aesencrypt.scala 200:36:@588.4]
  wire [7:0] _T_95; // @[aesencrypt.scala 201:18:@589.4]
  wire [7:0] _T_96; // @[aesencrypt.scala 245:27:@590.4]
  wire [7:0] _T_97; // @[aesencrypt.scala 245:34:@591.4]
  wire [7:0] _T_98; // @[aesencrypt.scala 249:22:@592.4]
  wire [8:0] _GEN_14; // @[aesencrypt.scala 198:27:@593.4]
  wire [8:0] _T_100; // @[aesencrypt.scala 198:27:@593.4]
  wire [8:0] _T_102; // @[aesencrypt.scala 198:35:@594.4]
  wire [7:0] _T_103; // @[aesencrypt.scala 198:46:@595.4]
  wire [7:0] _T_106; // @[aesencrypt.scala 199:31:@597.4]
  wire [7:0] _T_108; // @[aesencrypt.scala 200:25:@598.4]
  wire  _T_110; // @[aesencrypt.scala 200:36:@599.4]
  wire [7:0] _T_111; // @[aesencrypt.scala 201:18:@600.4]
  wire [7:0] _T_112; // @[aesencrypt.scala 251:23:@601.4]
  wire [7:0] _T_113; // @[aesencrypt.scala 251:30:@602.4]
  wire [7:0] _T_114; // @[aesencrypt.scala 254:25:@603.4]
  wire [8:0] _GEN_16; // @[aesencrypt.scala 198:27:@604.4]
  wire [8:0] _T_116; // @[aesencrypt.scala 198:27:@604.4]
  wire [8:0] _T_118; // @[aesencrypt.scala 198:35:@605.4]
  wire [7:0] _T_119; // @[aesencrypt.scala 198:46:@606.4]
  wire [7:0] _T_122; // @[aesencrypt.scala 199:31:@608.4]
  wire [7:0] _T_124; // @[aesencrypt.scala 200:25:@609.4]
  wire  _T_126; // @[aesencrypt.scala 200:36:@610.4]
  wire [7:0] _T_127; // @[aesencrypt.scala 201:18:@611.4]
  wire [7:0] _T_128; // @[aesencrypt.scala 256:25:@612.4]
  wire [7:0] _T_129; // @[aesencrypt.scala 256:32:@613.4]
  wire [15:0] _T_130; // @[Cat.scala 30:58:@614.4]
  wire [15:0] _T_131; // @[Cat.scala 30:58:@615.4]
  wire [31:0] _T_132; // @[Cat.scala 30:58:@616.4]
  wire [7:0] _T_133; // @[aesencrypt.scala 269:22:@617.4]
  wire [7:0] _T_134; // @[aesencrypt.scala 270:22:@618.4]
  wire [7:0] _T_135; // @[aesencrypt.scala 271:22:@619.4]
  wire [7:0] _T_136; // @[aesencrypt.scala 272:22:@620.4]
  wire [7:0] _T_137; // @[aesencrypt.scala 275:25:@621.4]
  wire [7:0] _T_138; // @[aesencrypt.scala 275:35:@622.4]
  wire [7:0] _T_139; // @[aesencrypt.scala 275:45:@623.4]
  wire [8:0] _GEN_18; // @[aesencrypt.scala 198:27:@625.4]
  wire [8:0] _T_142; // @[aesencrypt.scala 198:27:@625.4]
  wire [8:0] _T_144; // @[aesencrypt.scala 198:35:@626.4]
  wire [7:0] _T_145; // @[aesencrypt.scala 198:46:@627.4]
  wire [7:0] _T_148; // @[aesencrypt.scala 199:31:@629.4]
  wire [7:0] _T_150; // @[aesencrypt.scala 200:25:@630.4]
  wire  _T_152; // @[aesencrypt.scala 200:36:@631.4]
  wire [7:0] _T_153; // @[aesencrypt.scala 201:18:@632.4]
  wire [7:0] _T_154; // @[aesencrypt.scala 279:27:@633.4]
  wire [7:0] _T_155; // @[aesencrypt.scala 279:35:@634.4]
  wire [7:0] _T_156; // @[aesencrypt.scala 280:28:@635.4]
  wire [8:0] _GEN_20; // @[aesencrypt.scala 198:27:@636.4]
  wire [8:0] _T_158; // @[aesencrypt.scala 198:27:@636.4]
  wire [8:0] _T_160; // @[aesencrypt.scala 198:35:@637.4]
  wire [7:0] _T_161; // @[aesencrypt.scala 198:46:@638.4]
  wire [7:0] _T_164; // @[aesencrypt.scala 199:31:@640.4]
  wire [7:0] _T_166; // @[aesencrypt.scala 200:25:@641.4]
  wire  _T_168; // @[aesencrypt.scala 200:36:@642.4]
  wire [7:0] _T_169; // @[aesencrypt.scala 201:18:@643.4]
  wire [7:0] _T_170; // @[aesencrypt.scala 282:29:@644.4]
  wire [7:0] _T_171; // @[aesencrypt.scala 282:37:@645.4]
  wire [7:0] _T_172; // @[aesencrypt.scala 283:24:@646.4]
  wire [8:0] _GEN_22; // @[aesencrypt.scala 198:27:@647.4]
  wire [8:0] _T_174; // @[aesencrypt.scala 198:27:@647.4]
  wire [8:0] _T_176; // @[aesencrypt.scala 198:35:@648.4]
  wire [7:0] _T_177; // @[aesencrypt.scala 198:46:@649.4]
  wire [7:0] _T_180; // @[aesencrypt.scala 199:31:@651.4]
  wire [7:0] _T_182; // @[aesencrypt.scala 200:25:@652.4]
  wire  _T_184; // @[aesencrypt.scala 200:36:@653.4]
  wire [7:0] _T_185; // @[aesencrypt.scala 201:18:@654.4]
  wire [7:0] _T_186; // @[aesencrypt.scala 285:25:@655.4]
  wire [7:0] _T_187; // @[aesencrypt.scala 285:33:@656.4]
  wire [7:0] _T_188; // @[aesencrypt.scala 286:27:@657.4]
  wire [8:0] _GEN_24; // @[aesencrypt.scala 198:27:@658.4]
  wire [8:0] _T_190; // @[aesencrypt.scala 198:27:@658.4]
  wire [8:0] _T_192; // @[aesencrypt.scala 198:35:@659.4]
  wire [7:0] _T_193; // @[aesencrypt.scala 198:46:@660.4]
  wire [7:0] _T_196; // @[aesencrypt.scala 199:31:@662.4]
  wire [7:0] _T_198; // @[aesencrypt.scala 200:25:@663.4]
  wire  _T_200; // @[aesencrypt.scala 200:36:@664.4]
  wire [7:0] _T_201; // @[aesencrypt.scala 201:18:@665.4]
  wire [7:0] _T_202; // @[aesencrypt.scala 288:27:@666.4]
  wire [7:0] _T_203; // @[aesencrypt.scala 288:35:@667.4]
  wire [15:0] _T_204; // @[Cat.scala 30:58:@668.4]
  wire [15:0] _T_205; // @[Cat.scala 30:58:@669.4]
  wire [31:0] _T_206; // @[Cat.scala 30:58:@670.4]
  wire [7:0] _T_207; // @[aesencrypt.scala 301:26:@671.4]
  wire [7:0] _T_208; // @[aesencrypt.scala 302:26:@672.4]
  wire [7:0] _T_209; // @[aesencrypt.scala 303:26:@673.4]
  wire [7:0] _T_210; // @[aesencrypt.scala 304:26:@674.4]
  wire [7:0] _T_211; // @[aesencrypt.scala 307:25:@675.4]
  wire [7:0] _T_212; // @[aesencrypt.scala 307:35:@676.4]
  wire [7:0] _T_213; // @[aesencrypt.scala 307:45:@677.4]
  wire [8:0] _GEN_26; // @[aesencrypt.scala 198:27:@679.4]
  wire [8:0] _T_216; // @[aesencrypt.scala 198:27:@679.4]
  wire [8:0] _T_218; // @[aesencrypt.scala 198:35:@680.4]
  wire [7:0] _T_219; // @[aesencrypt.scala 198:46:@681.4]
  wire [7:0] _T_222; // @[aesencrypt.scala 199:31:@683.4]
  wire [7:0] _T_224; // @[aesencrypt.scala 200:25:@684.4]
  wire  _T_226; // @[aesencrypt.scala 200:36:@685.4]
  wire [7:0] _T_227; // @[aesencrypt.scala 201:18:@686.4]
  wire [7:0] _T_228; // @[aesencrypt.scala 311:27:@687.4]
  wire [7:0] _T_229; // @[aesencrypt.scala 311:35:@688.4]
  wire [7:0] _T_230; // @[aesencrypt.scala 312:28:@689.4]
  wire [8:0] _GEN_28; // @[aesencrypt.scala 198:27:@690.4]
  wire [8:0] _T_232; // @[aesencrypt.scala 198:27:@690.4]
  wire [8:0] _T_234; // @[aesencrypt.scala 198:35:@691.4]
  wire [7:0] _T_235; // @[aesencrypt.scala 198:46:@692.4]
  wire [7:0] _T_238; // @[aesencrypt.scala 199:31:@694.4]
  wire [7:0] _T_240; // @[aesencrypt.scala 200:25:@695.4]
  wire  _T_242; // @[aesencrypt.scala 200:36:@696.4]
  wire [7:0] _T_243; // @[aesencrypt.scala 201:18:@697.4]
  wire [7:0] _T_244; // @[aesencrypt.scala 314:29:@698.4]
  wire [7:0] _T_245; // @[aesencrypt.scala 314:37:@699.4]
  wire [7:0] _T_246; // @[aesencrypt.scala 315:24:@700.4]
  wire [8:0] _GEN_30; // @[aesencrypt.scala 198:27:@701.4]
  wire [8:0] _T_248; // @[aesencrypt.scala 198:27:@701.4]
  wire [8:0] _T_250; // @[aesencrypt.scala 198:35:@702.4]
  wire [7:0] _T_251; // @[aesencrypt.scala 198:46:@703.4]
  wire [7:0] _T_254; // @[aesencrypt.scala 199:31:@705.4]
  wire [7:0] _T_256; // @[aesencrypt.scala 200:25:@706.4]
  wire  _T_258; // @[aesencrypt.scala 200:36:@707.4]
  wire [7:0] _T_259; // @[aesencrypt.scala 201:18:@708.4]
  wire [7:0] _T_260; // @[aesencrypt.scala 317:25:@709.4]
  wire [7:0] _T_261; // @[aesencrypt.scala 317:33:@710.4]
  wire [7:0] _T_262; // @[aesencrypt.scala 318:27:@711.4]
  wire [8:0] _GEN_32; // @[aesencrypt.scala 198:27:@712.4]
  wire [8:0] _T_264; // @[aesencrypt.scala 198:27:@712.4]
  wire [8:0] _T_266; // @[aesencrypt.scala 198:35:@713.4]
  wire [7:0] _T_267; // @[aesencrypt.scala 198:46:@714.4]
  wire [7:0] _T_270; // @[aesencrypt.scala 199:31:@716.4]
  wire [7:0] _T_272; // @[aesencrypt.scala 200:25:@717.4]
  wire  _T_274; // @[aesencrypt.scala 200:36:@718.4]
  wire [7:0] _T_275; // @[aesencrypt.scala 201:18:@719.4]
  wire [7:0] _T_276; // @[aesencrypt.scala 320:27:@720.4]
  wire [7:0] _T_277; // @[aesencrypt.scala 320:35:@721.4]
  wire [15:0] _T_278; // @[Cat.scala 30:58:@722.4]
  wire [15:0] _T_279; // @[Cat.scala 30:58:@723.4]
  wire [31:0] _T_280; // @[Cat.scala 30:58:@724.4]
  wire [7:0] _T_281; // @[aesencrypt.scala 333:22:@725.4]
  wire [7:0] _T_282; // @[aesencrypt.scala 334:22:@726.4]
  wire [7:0] _T_283; // @[aesencrypt.scala 335:22:@727.4]
  wire [7:0] _T_284; // @[aesencrypt.scala 336:22:@728.4]
  wire [7:0] _T_285; // @[aesencrypt.scala 340:25:@729.4]
  wire [7:0] _T_286; // @[aesencrypt.scala 340:35:@730.4]
  wire [7:0] _T_287; // @[aesencrypt.scala 340:45:@731.4]
  wire [8:0] _GEN_34; // @[aesencrypt.scala 198:27:@733.4]
  wire [8:0] _T_290; // @[aesencrypt.scala 198:27:@733.4]
  wire [8:0] _T_292; // @[aesencrypt.scala 198:35:@734.4]
  wire [7:0] _T_293; // @[aesencrypt.scala 198:46:@735.4]
  wire [7:0] _T_296; // @[aesencrypt.scala 199:31:@737.4]
  wire [7:0] _T_298; // @[aesencrypt.scala 200:25:@738.4]
  wire  _T_300; // @[aesencrypt.scala 200:36:@739.4]
  wire [7:0] _T_301; // @[aesencrypt.scala 201:18:@740.4]
  wire [7:0] _T_302; // @[aesencrypt.scala 344:27:@741.4]
  wire [7:0] _T_303; // @[aesencrypt.scala 344:35:@742.4]
  wire [7:0] _T_304; // @[aesencrypt.scala 345:28:@743.4]
  wire [8:0] _GEN_36; // @[aesencrypt.scala 198:27:@744.4]
  wire [8:0] _T_306; // @[aesencrypt.scala 198:27:@744.4]
  wire [8:0] _T_308; // @[aesencrypt.scala 198:35:@745.4]
  wire [7:0] _T_309; // @[aesencrypt.scala 198:46:@746.4]
  wire [7:0] _T_312; // @[aesencrypt.scala 199:31:@748.4]
  wire [7:0] _T_314; // @[aesencrypt.scala 200:25:@749.4]
  wire  _T_316; // @[aesencrypt.scala 200:36:@750.4]
  wire [7:0] _T_317; // @[aesencrypt.scala 201:18:@751.4]
  wire [7:0] _T_318; // @[aesencrypt.scala 347:29:@752.4]
  wire [7:0] _T_319; // @[aesencrypt.scala 347:37:@753.4]
  wire [7:0] _T_320; // @[aesencrypt.scala 348:24:@754.4]
  wire [8:0] _GEN_38; // @[aesencrypt.scala 198:27:@755.4]
  wire [8:0] _T_322; // @[aesencrypt.scala 198:27:@755.4]
  wire [8:0] _T_324; // @[aesencrypt.scala 198:35:@756.4]
  wire [7:0] _T_325; // @[aesencrypt.scala 198:46:@757.4]
  wire [7:0] _T_328; // @[aesencrypt.scala 199:31:@759.4]
  wire [7:0] _T_330; // @[aesencrypt.scala 200:25:@760.4]
  wire  _T_332; // @[aesencrypt.scala 200:36:@761.4]
  wire [7:0] _T_333; // @[aesencrypt.scala 201:18:@762.4]
  wire [7:0] _T_334; // @[aesencrypt.scala 350:25:@763.4]
  wire [7:0] _T_335; // @[aesencrypt.scala 350:33:@764.4]
  wire [7:0] _T_336; // @[aesencrypt.scala 351:27:@765.4]
  wire [8:0] _GEN_40; // @[aesencrypt.scala 198:27:@766.4]
  wire [8:0] _T_338; // @[aesencrypt.scala 198:27:@766.4]
  wire [8:0] _T_340; // @[aesencrypt.scala 198:35:@767.4]
  wire [7:0] _T_341; // @[aesencrypt.scala 198:46:@768.4]
  wire [7:0] _T_344; // @[aesencrypt.scala 199:31:@770.4]
  wire [7:0] _T_346; // @[aesencrypt.scala 200:25:@771.4]
  wire  _T_348; // @[aesencrypt.scala 200:36:@772.4]
  wire [7:0] _T_349; // @[aesencrypt.scala 201:18:@773.4]
  wire [7:0] _T_350; // @[aesencrypt.scala 353:27:@774.4]
  wire [7:0] _T_351; // @[aesencrypt.scala 353:35:@775.4]
  wire [15:0] _T_352; // @[Cat.scala 30:58:@776.4]
  wire [15:0] _T_353; // @[Cat.scala 30:58:@777.4]
  wire [31:0] _T_354; // @[Cat.scala 30:58:@778.4]
  wire [63:0] _T_355; // @[Cat.scala 30:58:@779.4]
  wire [63:0] _T_356; // @[Cat.scala 30:58:@780.4]
  wire [127:0] state2; // @[Cat.scala 30:58:@781.4]
  wire [127:0] state3; // @[aesencrypt.scala 156:25:@782.4]
  wire [127:0] state31; // @[aesencrypt.scala 156:25:@815.4]
  wire  _T_389; // @[Mux.scala 46:19:@817.4]
  wire [127:0] _T_390; // @[Mux.scala 46:16:@818.4]
  wire  _T_391; // @[Mux.scala 46:19:@819.4]
  wire [127:0] output$; // @[Mux.scala 46:16:@820.4]
  wire [127:0] _T_394; // @[aesencrypt.scala 74:16:@822.4]
  wire  _T_396; // @[aesencrypt.scala 84:27:@826.8]
  wire  _T_398; // @[aesencrypt.scala 97:33:@831.10]
  wire  _T_400; // @[aesencrypt.scala 97:55:@832.10]
  wire  _T_401; // @[aesencrypt.scala 97:39:@833.10]
  wire [3:0] _GEN_0; // @[aesencrypt.scala 124:9:@839.12]
  wire [127:0] _GEN_2; // @[aesencrypt.scala 97:63:@834.10]
  wire [3:0] _GEN_3; // @[aesencrypt.scala 97:63:@834.10]
  wire [127:0] _GEN_4; // @[aesencrypt.scala 85:9:@827.8]
  wire [3:0] _GEN_5; // @[aesencrypt.scala 85:9:@827.8]
  wire [127:0] _GEN_8; // @[aesencrypt.scala 78:3:@824.4]
  wire [3:0] _GEN_9; // @[aesencrypt.scala 78:3:@824.4]
  assign _T_19 = roundCounter == 4'ha; // @[aesencrypt.scala 24:37:@521.4]
  assign _T_21 = io_en ? _T_19 : 1'h0; // @[aesencrypt.scala 24:17:@522.4]
  assign _T_23 = roundCounter + 4'h1; // @[aesencrypt.scala 43:42:@524.4]
  assign _T_24 = _T_23[3:0]; // @[aesencrypt.scala 43:42:@525.4]
  assign _T_26 = io_en ? _T_24 : 4'h0; // @[aesencrypt.scala 43:22:@526.4]
  assign _T_28 = io_en ? roundCounter : 4'h0; // @[aesencrypt.scala 44:21:@528.4]
  assign t = io_data ^ io_rkey; // @[aesencrypt.scala 156:25:@530.4]
  assign _T_29 = io_sio_data2[31:24]; // @[aesencrypt.scala 168:14:@532.4]
  assign _T_30 = io_sio_data2[119:112]; // @[aesencrypt.scala 169:14:@533.4]
  assign _T_31 = io_sio_data2[79:72]; // @[aesencrypt.scala 170:14:@534.4]
  assign _T_32 = io_sio_data2[39:32]; // @[aesencrypt.scala 171:14:@535.4]
  assign _T_33 = {_T_31,_T_32}; // @[Cat.scala 30:58:@536.4]
  assign _T_34 = {_T_29,_T_30}; // @[Cat.scala 30:58:@537.4]
  assign _T_35 = {_T_34,_T_33}; // @[Cat.scala 30:58:@538.4]
  assign _T_36 = io_sio_data2[63:56]; // @[aesencrypt.scala 174:15:@539.4]
  assign _T_37 = io_sio_data2[23:16]; // @[aesencrypt.scala 175:15:@540.4]
  assign _T_38 = io_sio_data2[111:104]; // @[aesencrypt.scala 177:14:@541.4]
  assign _T_39 = io_sio_data2[71:64]; // @[aesencrypt.scala 178:14:@542.4]
  assign _T_40 = {_T_38,_T_39}; // @[Cat.scala 30:58:@543.4]
  assign _T_41 = {_T_36,_T_37}; // @[Cat.scala 30:58:@544.4]
  assign _T_42 = {_T_41,_T_40}; // @[Cat.scala 30:58:@545.4]
  assign _T_43 = io_sio_data2[95:88]; // @[aesencrypt.scala 181:15:@546.4]
  assign _T_44 = io_sio_data2[55:48]; // @[aesencrypt.scala 182:15:@547.4]
  assign _T_45 = io_sio_data2[15:8]; // @[aesencrypt.scala 183:15:@548.4]
  assign _T_46 = io_sio_data2[103:96]; // @[aesencrypt.scala 184:15:@549.4]
  assign _T_47 = {_T_45,_T_46}; // @[Cat.scala 30:58:@550.4]
  assign _T_48 = {_T_43,_T_44}; // @[Cat.scala 30:58:@551.4]
  assign _T_49 = {_T_48,_T_47}; // @[Cat.scala 30:58:@552.4]
  assign _T_50 = io_sio_data2[127:120]; // @[aesencrypt.scala 187:14:@553.4]
  assign _T_51 = io_sio_data2[87:80]; // @[aesencrypt.scala 188:14:@554.4]
  assign _T_52 = io_sio_data2[47:40]; // @[aesencrypt.scala 189:14:@555.4]
  assign _T_53 = io_sio_data2[7:0]; // @[aesencrypt.scala 190:14:@556.4]
  assign _T_54 = {_T_52,_T_53}; // @[Cat.scala 30:58:@557.4]
  assign _T_55 = {_T_50,_T_51}; // @[Cat.scala 30:58:@558.4]
  assign _T_56 = {_T_55,_T_54}; // @[Cat.scala 30:58:@559.4]
  assign _T_57 = {_T_42,_T_35}; // @[Cat.scala 30:58:@560.4]
  assign _T_58 = {_T_56,_T_49}; // @[Cat.scala 30:58:@561.4]
  assign state1 = {_T_58,_T_57}; // @[Cat.scala 30:58:@562.4]
  assign _T_59 = state1[103:96]; // @[aesencrypt.scala 220:21:@563.4]
  assign _T_60 = state1[111:104]; // @[aesencrypt.scala 221:21:@564.4]
  assign _T_61 = state1[119:112]; // @[aesencrypt.scala 222:21:@565.4]
  assign _T_62 = state1[127:120]; // @[aesencrypt.scala 223:21:@566.4]
  assign _T_63 = _T_62 ^ _T_61; // @[aesencrypt.scala 231:23:@567.4]
  assign _T_64 = _T_63 ^ _T_60; // @[aesencrypt.scala 231:32:@568.4]
  assign _T_65 = _T_64 ^ _T_59; // @[aesencrypt.scala 231:41:@569.4]
  assign _GEN_10 = {{1'd0}, _T_63}; // @[aesencrypt.scala 198:27:@571.4]
  assign _T_68 = _GEN_10 << 1'h1; // @[aesencrypt.scala 198:27:@571.4]
  assign _T_70 = _T_68 ^ 9'h1b; // @[aesencrypt.scala 198:35:@572.4]
  assign _T_71 = _T_70[7:0]; // @[aesencrypt.scala 198:46:@573.4]
  assign _T_74 = _T_68[7:0]; // @[aesencrypt.scala 199:31:@575.4]
  assign _T_76 = _T_63 & 8'h80; // @[aesencrypt.scala 200:25:@576.4]
  assign _T_78 = _T_76 == 8'h80; // @[aesencrypt.scala 200:36:@577.4]
  assign _T_79 = _T_78 ? _T_71 : _T_74; // @[aesencrypt.scala 201:18:@578.4]
  assign _T_80 = _T_62 ^ _T_79; // @[aesencrypt.scala 238:25:@579.4]
  assign _T_81 = _T_80 ^ _T_65; // @[aesencrypt.scala 238:32:@580.4]
  assign _T_82 = _T_61 ^ _T_60; // @[aesencrypt.scala 241:26:@581.4]
  assign _GEN_12 = {{1'd0}, _T_82}; // @[aesencrypt.scala 198:27:@582.4]
  assign _T_84 = _GEN_12 << 1'h1; // @[aesencrypt.scala 198:27:@582.4]
  assign _T_86 = _T_84 ^ 9'h1b; // @[aesencrypt.scala 198:35:@583.4]
  assign _T_87 = _T_86[7:0]; // @[aesencrypt.scala 198:46:@584.4]
  assign _T_90 = _T_84[7:0]; // @[aesencrypt.scala 199:31:@586.4]
  assign _T_92 = _T_82 & 8'h80; // @[aesencrypt.scala 200:25:@587.4]
  assign _T_94 = _T_92 == 8'h80; // @[aesencrypt.scala 200:36:@588.4]
  assign _T_95 = _T_94 ? _T_87 : _T_90; // @[aesencrypt.scala 201:18:@589.4]
  assign _T_96 = _T_61 ^ _T_95; // @[aesencrypt.scala 245:27:@590.4]
  assign _T_97 = _T_96 ^ _T_65; // @[aesencrypt.scala 245:34:@591.4]
  assign _T_98 = _T_60 ^ _T_59; // @[aesencrypt.scala 249:22:@592.4]
  assign _GEN_14 = {{1'd0}, _T_98}; // @[aesencrypt.scala 198:27:@593.4]
  assign _T_100 = _GEN_14 << 1'h1; // @[aesencrypt.scala 198:27:@593.4]
  assign _T_102 = _T_100 ^ 9'h1b; // @[aesencrypt.scala 198:35:@594.4]
  assign _T_103 = _T_102[7:0]; // @[aesencrypt.scala 198:46:@595.4]
  assign _T_106 = _T_100[7:0]; // @[aesencrypt.scala 199:31:@597.4]
  assign _T_108 = _T_98 & 8'h80; // @[aesencrypt.scala 200:25:@598.4]
  assign _T_110 = _T_108 == 8'h80; // @[aesencrypt.scala 200:36:@599.4]
  assign _T_111 = _T_110 ? _T_103 : _T_106; // @[aesencrypt.scala 201:18:@600.4]
  assign _T_112 = _T_60 ^ _T_111; // @[aesencrypt.scala 251:23:@601.4]
  assign _T_113 = _T_112 ^ _T_65; // @[aesencrypt.scala 251:30:@602.4]
  assign _T_114 = _T_59 ^ _T_62; // @[aesencrypt.scala 254:25:@603.4]
  assign _GEN_16 = {{1'd0}, _T_114}; // @[aesencrypt.scala 198:27:@604.4]
  assign _T_116 = _GEN_16 << 1'h1; // @[aesencrypt.scala 198:27:@604.4]
  assign _T_118 = _T_116 ^ 9'h1b; // @[aesencrypt.scala 198:35:@605.4]
  assign _T_119 = _T_118[7:0]; // @[aesencrypt.scala 198:46:@606.4]
  assign _T_122 = _T_116[7:0]; // @[aesencrypt.scala 199:31:@608.4]
  assign _T_124 = _T_114 & 8'h80; // @[aesencrypt.scala 200:25:@609.4]
  assign _T_126 = _T_124 == 8'h80; // @[aesencrypt.scala 200:36:@610.4]
  assign _T_127 = _T_126 ? _T_119 : _T_122; // @[aesencrypt.scala 201:18:@611.4]
  assign _T_128 = _T_59 ^ _T_127; // @[aesencrypt.scala 256:25:@612.4]
  assign _T_129 = _T_128 ^ _T_65; // @[aesencrypt.scala 256:32:@613.4]
  assign _T_130 = {_T_113,_T_129}; // @[Cat.scala 30:58:@614.4]
  assign _T_131 = {_T_81,_T_97}; // @[Cat.scala 30:58:@615.4]
  assign _T_132 = {_T_131,_T_130}; // @[Cat.scala 30:58:@616.4]
  assign _T_133 = state1[71:64]; // @[aesencrypt.scala 269:22:@617.4]
  assign _T_134 = state1[79:72]; // @[aesencrypt.scala 270:22:@618.4]
  assign _T_135 = state1[87:80]; // @[aesencrypt.scala 271:22:@619.4]
  assign _T_136 = state1[95:88]; // @[aesencrypt.scala 272:22:@620.4]
  assign _T_137 = _T_136 ^ _T_135; // @[aesencrypt.scala 275:25:@621.4]
  assign _T_138 = _T_137 ^ _T_134; // @[aesencrypt.scala 275:35:@622.4]
  assign _T_139 = _T_138 ^ _T_133; // @[aesencrypt.scala 275:45:@623.4]
  assign _GEN_18 = {{1'd0}, _T_137}; // @[aesencrypt.scala 198:27:@625.4]
  assign _T_142 = _GEN_18 << 1'h1; // @[aesencrypt.scala 198:27:@625.4]
  assign _T_144 = _T_142 ^ 9'h1b; // @[aesencrypt.scala 198:35:@626.4]
  assign _T_145 = _T_144[7:0]; // @[aesencrypt.scala 198:46:@627.4]
  assign _T_148 = _T_142[7:0]; // @[aesencrypt.scala 199:31:@629.4]
  assign _T_150 = _T_137 & 8'h80; // @[aesencrypt.scala 200:25:@630.4]
  assign _T_152 = _T_150 == 8'h80; // @[aesencrypt.scala 200:36:@631.4]
  assign _T_153 = _T_152 ? _T_145 : _T_148; // @[aesencrypt.scala 201:18:@632.4]
  assign _T_154 = _T_136 ^ _T_153; // @[aesencrypt.scala 279:27:@633.4]
  assign _T_155 = _T_154 ^ _T_139; // @[aesencrypt.scala 279:35:@634.4]
  assign _T_156 = _T_135 ^ _T_134; // @[aesencrypt.scala 280:28:@635.4]
  assign _GEN_20 = {{1'd0}, _T_156}; // @[aesencrypt.scala 198:27:@636.4]
  assign _T_158 = _GEN_20 << 1'h1; // @[aesencrypt.scala 198:27:@636.4]
  assign _T_160 = _T_158 ^ 9'h1b; // @[aesencrypt.scala 198:35:@637.4]
  assign _T_161 = _T_160[7:0]; // @[aesencrypt.scala 198:46:@638.4]
  assign _T_164 = _T_158[7:0]; // @[aesencrypt.scala 199:31:@640.4]
  assign _T_166 = _T_156 & 8'h80; // @[aesencrypt.scala 200:25:@641.4]
  assign _T_168 = _T_166 == 8'h80; // @[aesencrypt.scala 200:36:@642.4]
  assign _T_169 = _T_168 ? _T_161 : _T_164; // @[aesencrypt.scala 201:18:@643.4]
  assign _T_170 = _T_135 ^ _T_169; // @[aesencrypt.scala 282:29:@644.4]
  assign _T_171 = _T_170 ^ _T_139; // @[aesencrypt.scala 282:37:@645.4]
  assign _T_172 = _T_134 ^ _T_133; // @[aesencrypt.scala 283:24:@646.4]
  assign _GEN_22 = {{1'd0}, _T_172}; // @[aesencrypt.scala 198:27:@647.4]
  assign _T_174 = _GEN_22 << 1'h1; // @[aesencrypt.scala 198:27:@647.4]
  assign _T_176 = _T_174 ^ 9'h1b; // @[aesencrypt.scala 198:35:@648.4]
  assign _T_177 = _T_176[7:0]; // @[aesencrypt.scala 198:46:@649.4]
  assign _T_180 = _T_174[7:0]; // @[aesencrypt.scala 199:31:@651.4]
  assign _T_182 = _T_172 & 8'h80; // @[aesencrypt.scala 200:25:@652.4]
  assign _T_184 = _T_182 == 8'h80; // @[aesencrypt.scala 200:36:@653.4]
  assign _T_185 = _T_184 ? _T_177 : _T_180; // @[aesencrypt.scala 201:18:@654.4]
  assign _T_186 = _T_134 ^ _T_185; // @[aesencrypt.scala 285:25:@655.4]
  assign _T_187 = _T_186 ^ _T_139; // @[aesencrypt.scala 285:33:@656.4]
  assign _T_188 = _T_133 ^ _T_136; // @[aesencrypt.scala 286:27:@657.4]
  assign _GEN_24 = {{1'd0}, _T_188}; // @[aesencrypt.scala 198:27:@658.4]
  assign _T_190 = _GEN_24 << 1'h1; // @[aesencrypt.scala 198:27:@658.4]
  assign _T_192 = _T_190 ^ 9'h1b; // @[aesencrypt.scala 198:35:@659.4]
  assign _T_193 = _T_192[7:0]; // @[aesencrypt.scala 198:46:@660.4]
  assign _T_196 = _T_190[7:0]; // @[aesencrypt.scala 199:31:@662.4]
  assign _T_198 = _T_188 & 8'h80; // @[aesencrypt.scala 200:25:@663.4]
  assign _T_200 = _T_198 == 8'h80; // @[aesencrypt.scala 200:36:@664.4]
  assign _T_201 = _T_200 ? _T_193 : _T_196; // @[aesencrypt.scala 201:18:@665.4]
  assign _T_202 = _T_133 ^ _T_201; // @[aesencrypt.scala 288:27:@666.4]
  assign _T_203 = _T_202 ^ _T_139; // @[aesencrypt.scala 288:35:@667.4]
  assign _T_204 = {_T_187,_T_203}; // @[Cat.scala 30:58:@668.4]
  assign _T_205 = {_T_155,_T_171}; // @[Cat.scala 30:58:@669.4]
  assign _T_206 = {_T_205,_T_204}; // @[Cat.scala 30:58:@670.4]
  assign _T_207 = state1[39:32]; // @[aesencrypt.scala 301:26:@671.4]
  assign _T_208 = state1[47:40]; // @[aesencrypt.scala 302:26:@672.4]
  assign _T_209 = state1[55:48]; // @[aesencrypt.scala 303:26:@673.4]
  assign _T_210 = state1[63:56]; // @[aesencrypt.scala 304:26:@674.4]
  assign _T_211 = _T_210 ^ _T_209; // @[aesencrypt.scala 307:25:@675.4]
  assign _T_212 = _T_211 ^ _T_208; // @[aesencrypt.scala 307:35:@676.4]
  assign _T_213 = _T_212 ^ _T_207; // @[aesencrypt.scala 307:45:@677.4]
  assign _GEN_26 = {{1'd0}, _T_211}; // @[aesencrypt.scala 198:27:@679.4]
  assign _T_216 = _GEN_26 << 1'h1; // @[aesencrypt.scala 198:27:@679.4]
  assign _T_218 = _T_216 ^ 9'h1b; // @[aesencrypt.scala 198:35:@680.4]
  assign _T_219 = _T_218[7:0]; // @[aesencrypt.scala 198:46:@681.4]
  assign _T_222 = _T_216[7:0]; // @[aesencrypt.scala 199:31:@683.4]
  assign _T_224 = _T_211 & 8'h80; // @[aesencrypt.scala 200:25:@684.4]
  assign _T_226 = _T_224 == 8'h80; // @[aesencrypt.scala 200:36:@685.4]
  assign _T_227 = _T_226 ? _T_219 : _T_222; // @[aesencrypt.scala 201:18:@686.4]
  assign _T_228 = _T_210 ^ _T_227; // @[aesencrypt.scala 311:27:@687.4]
  assign _T_229 = _T_228 ^ _T_213; // @[aesencrypt.scala 311:35:@688.4]
  assign _T_230 = _T_209 ^ _T_208; // @[aesencrypt.scala 312:28:@689.4]
  assign _GEN_28 = {{1'd0}, _T_230}; // @[aesencrypt.scala 198:27:@690.4]
  assign _T_232 = _GEN_28 << 1'h1; // @[aesencrypt.scala 198:27:@690.4]
  assign _T_234 = _T_232 ^ 9'h1b; // @[aesencrypt.scala 198:35:@691.4]
  assign _T_235 = _T_234[7:0]; // @[aesencrypt.scala 198:46:@692.4]
  assign _T_238 = _T_232[7:0]; // @[aesencrypt.scala 199:31:@694.4]
  assign _T_240 = _T_230 & 8'h80; // @[aesencrypt.scala 200:25:@695.4]
  assign _T_242 = _T_240 == 8'h80; // @[aesencrypt.scala 200:36:@696.4]
  assign _T_243 = _T_242 ? _T_235 : _T_238; // @[aesencrypt.scala 201:18:@697.4]
  assign _T_244 = _T_209 ^ _T_243; // @[aesencrypt.scala 314:29:@698.4]
  assign _T_245 = _T_244 ^ _T_213; // @[aesencrypt.scala 314:37:@699.4]
  assign _T_246 = _T_208 ^ _T_207; // @[aesencrypt.scala 315:24:@700.4]
  assign _GEN_30 = {{1'd0}, _T_246}; // @[aesencrypt.scala 198:27:@701.4]
  assign _T_248 = _GEN_30 << 1'h1; // @[aesencrypt.scala 198:27:@701.4]
  assign _T_250 = _T_248 ^ 9'h1b; // @[aesencrypt.scala 198:35:@702.4]
  assign _T_251 = _T_250[7:0]; // @[aesencrypt.scala 198:46:@703.4]
  assign _T_254 = _T_248[7:0]; // @[aesencrypt.scala 199:31:@705.4]
  assign _T_256 = _T_246 & 8'h80; // @[aesencrypt.scala 200:25:@706.4]
  assign _T_258 = _T_256 == 8'h80; // @[aesencrypt.scala 200:36:@707.4]
  assign _T_259 = _T_258 ? _T_251 : _T_254; // @[aesencrypt.scala 201:18:@708.4]
  assign _T_260 = _T_208 ^ _T_259; // @[aesencrypt.scala 317:25:@709.4]
  assign _T_261 = _T_260 ^ _T_213; // @[aesencrypt.scala 317:33:@710.4]
  assign _T_262 = _T_207 ^ _T_210; // @[aesencrypt.scala 318:27:@711.4]
  assign _GEN_32 = {{1'd0}, _T_262}; // @[aesencrypt.scala 198:27:@712.4]
  assign _T_264 = _GEN_32 << 1'h1; // @[aesencrypt.scala 198:27:@712.4]
  assign _T_266 = _T_264 ^ 9'h1b; // @[aesencrypt.scala 198:35:@713.4]
  assign _T_267 = _T_266[7:0]; // @[aesencrypt.scala 198:46:@714.4]
  assign _T_270 = _T_264[7:0]; // @[aesencrypt.scala 199:31:@716.4]
  assign _T_272 = _T_262 & 8'h80; // @[aesencrypt.scala 200:25:@717.4]
  assign _T_274 = _T_272 == 8'h80; // @[aesencrypt.scala 200:36:@718.4]
  assign _T_275 = _T_274 ? _T_267 : _T_270; // @[aesencrypt.scala 201:18:@719.4]
  assign _T_276 = _T_207 ^ _T_275; // @[aesencrypt.scala 320:27:@720.4]
  assign _T_277 = _T_276 ^ _T_213; // @[aesencrypt.scala 320:35:@721.4]
  assign _T_278 = {_T_261,_T_277}; // @[Cat.scala 30:58:@722.4]
  assign _T_279 = {_T_229,_T_245}; // @[Cat.scala 30:58:@723.4]
  assign _T_280 = {_T_279,_T_278}; // @[Cat.scala 30:58:@724.4]
  assign _T_281 = state1[7:0]; // @[aesencrypt.scala 333:22:@725.4]
  assign _T_282 = state1[15:8]; // @[aesencrypt.scala 334:22:@726.4]
  assign _T_283 = state1[23:16]; // @[aesencrypt.scala 335:22:@727.4]
  assign _T_284 = state1[31:24]; // @[aesencrypt.scala 336:22:@728.4]
  assign _T_285 = _T_284 ^ _T_283; // @[aesencrypt.scala 340:25:@729.4]
  assign _T_286 = _T_285 ^ _T_282; // @[aesencrypt.scala 340:35:@730.4]
  assign _T_287 = _T_286 ^ _T_281; // @[aesencrypt.scala 340:45:@731.4]
  assign _GEN_34 = {{1'd0}, _T_285}; // @[aesencrypt.scala 198:27:@733.4]
  assign _T_290 = _GEN_34 << 1'h1; // @[aesencrypt.scala 198:27:@733.4]
  assign _T_292 = _T_290 ^ 9'h1b; // @[aesencrypt.scala 198:35:@734.4]
  assign _T_293 = _T_292[7:0]; // @[aesencrypt.scala 198:46:@735.4]
  assign _T_296 = _T_290[7:0]; // @[aesencrypt.scala 199:31:@737.4]
  assign _T_298 = _T_285 & 8'h80; // @[aesencrypt.scala 200:25:@738.4]
  assign _T_300 = _T_298 == 8'h80; // @[aesencrypt.scala 200:36:@739.4]
  assign _T_301 = _T_300 ? _T_293 : _T_296; // @[aesencrypt.scala 201:18:@740.4]
  assign _T_302 = _T_284 ^ _T_301; // @[aesencrypt.scala 344:27:@741.4]
  assign _T_303 = _T_302 ^ _T_287; // @[aesencrypt.scala 344:35:@742.4]
  assign _T_304 = _T_283 ^ _T_282; // @[aesencrypt.scala 345:28:@743.4]
  assign _GEN_36 = {{1'd0}, _T_304}; // @[aesencrypt.scala 198:27:@744.4]
  assign _T_306 = _GEN_36 << 1'h1; // @[aesencrypt.scala 198:27:@744.4]
  assign _T_308 = _T_306 ^ 9'h1b; // @[aesencrypt.scala 198:35:@745.4]
  assign _T_309 = _T_308[7:0]; // @[aesencrypt.scala 198:46:@746.4]
  assign _T_312 = _T_306[7:0]; // @[aesencrypt.scala 199:31:@748.4]
  assign _T_314 = _T_304 & 8'h80; // @[aesencrypt.scala 200:25:@749.4]
  assign _T_316 = _T_314 == 8'h80; // @[aesencrypt.scala 200:36:@750.4]
  assign _T_317 = _T_316 ? _T_309 : _T_312; // @[aesencrypt.scala 201:18:@751.4]
  assign _T_318 = _T_283 ^ _T_317; // @[aesencrypt.scala 347:29:@752.4]
  assign _T_319 = _T_318 ^ _T_287; // @[aesencrypt.scala 347:37:@753.4]
  assign _T_320 = _T_282 ^ _T_281; // @[aesencrypt.scala 348:24:@754.4]
  assign _GEN_38 = {{1'd0}, _T_320}; // @[aesencrypt.scala 198:27:@755.4]
  assign _T_322 = _GEN_38 << 1'h1; // @[aesencrypt.scala 198:27:@755.4]
  assign _T_324 = _T_322 ^ 9'h1b; // @[aesencrypt.scala 198:35:@756.4]
  assign _T_325 = _T_324[7:0]; // @[aesencrypt.scala 198:46:@757.4]
  assign _T_328 = _T_322[7:0]; // @[aesencrypt.scala 199:31:@759.4]
  assign _T_330 = _T_320 & 8'h80; // @[aesencrypt.scala 200:25:@760.4]
  assign _T_332 = _T_330 == 8'h80; // @[aesencrypt.scala 200:36:@761.4]
  assign _T_333 = _T_332 ? _T_325 : _T_328; // @[aesencrypt.scala 201:18:@762.4]
  assign _T_334 = _T_282 ^ _T_333; // @[aesencrypt.scala 350:25:@763.4]
  assign _T_335 = _T_334 ^ _T_287; // @[aesencrypt.scala 350:33:@764.4]
  assign _T_336 = _T_281 ^ _T_284; // @[aesencrypt.scala 351:27:@765.4]
  assign _GEN_40 = {{1'd0}, _T_336}; // @[aesencrypt.scala 198:27:@766.4]
  assign _T_338 = _GEN_40 << 1'h1; // @[aesencrypt.scala 198:27:@766.4]
  assign _T_340 = _T_338 ^ 9'h1b; // @[aesencrypt.scala 198:35:@767.4]
  assign _T_341 = _T_340[7:0]; // @[aesencrypt.scala 198:46:@768.4]
  assign _T_344 = _T_338[7:0]; // @[aesencrypt.scala 199:31:@770.4]
  assign _T_346 = _T_336 & 8'h80; // @[aesencrypt.scala 200:25:@771.4]
  assign _T_348 = _T_346 == 8'h80; // @[aesencrypt.scala 200:36:@772.4]
  assign _T_349 = _T_348 ? _T_341 : _T_344; // @[aesencrypt.scala 201:18:@773.4]
  assign _T_350 = _T_281 ^ _T_349; // @[aesencrypt.scala 353:27:@774.4]
  assign _T_351 = _T_350 ^ _T_287; // @[aesencrypt.scala 353:35:@775.4]
  assign _T_352 = {_T_335,_T_351}; // @[Cat.scala 30:58:@776.4]
  assign _T_353 = {_T_303,_T_319}; // @[Cat.scala 30:58:@777.4]
  assign _T_354 = {_T_353,_T_352}; // @[Cat.scala 30:58:@778.4]
  assign _T_355 = {_T_280,_T_354}; // @[Cat.scala 30:58:@779.4]
  assign _T_356 = {_T_132,_T_206}; // @[Cat.scala 30:58:@780.4]
  assign state2 = {_T_356,_T_355}; // @[Cat.scala 30:58:@781.4]
  assign state3 = state2 ^ io_rkey; // @[aesencrypt.scala 156:25:@782.4]
  assign state31 = state1 ^ io_rkey; // @[aesencrypt.scala 156:25:@815.4]
  assign _T_389 = 4'ha == roundCounter; // @[Mux.scala 46:19:@817.4]
  assign _T_390 = _T_389 ? state31 : state3; // @[Mux.scala 46:16:@818.4]
  assign _T_391 = 4'h0 == roundCounter; // @[Mux.scala 46:19:@819.4]
  assign output$ = _T_391 ? t : _T_390; // @[Mux.scala 46:16:@820.4]
  assign _T_394 = io_en ? output$ : 128'h0; // @[aesencrypt.scala 74:16:@822.4]
  assign _T_396 = roundCounter == 4'h0; // @[aesencrypt.scala 84:27:@826.8]
  assign _T_398 = roundCounter > 4'h0; // @[aesencrypt.scala 97:33:@831.10]
  assign _T_400 = roundCounter <= 4'h9; // @[aesencrypt.scala 97:55:@832.10]
  assign _T_401 = _T_398 & _T_400; // @[aesencrypt.scala 97:39:@833.10]
  assign _GEN_0 = _T_19 ? 4'h0 : _T_26; // @[aesencrypt.scala 124:9:@839.12]
  assign _GEN_2 = _T_401 ? state3 : state31; // @[aesencrypt.scala 97:63:@834.10]
  assign _GEN_3 = _T_401 ? _T_26 : _GEN_0; // @[aesencrypt.scala 97:63:@834.10]
  assign _GEN_4 = _T_396 ? t : _GEN_2; // @[aesencrypt.scala 85:9:@827.8]
  assign _GEN_5 = _T_396 ? _T_26 : _GEN_3; // @[aesencrypt.scala 85:9:@827.8]
  assign _GEN_8 = io_en ? _GEN_4 : state31; // @[aesencrypt.scala 78:3:@824.4]
  assign _GEN_9 = io_en ? _GEN_5 : _T_26; // @[aesencrypt.scala 78:3:@824.4]
  assign io_done = _T_21;
  assign io_sio_addr2 = state;
  assign io_out = _T_394;
  assign io_roundOut = _T_28;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  roundCounter = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{$random}};
  state = _RAND_1[127:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      roundCounter <= 4'hf;
    end else begin
      if (io_en) begin
        if (_T_396) begin
          if (io_en) begin
            roundCounter <= _T_24;
          end else begin
            roundCounter <= 4'h0;
          end
        end else begin
          if (_T_401) begin
            if (io_en) begin
              roundCounter <= _T_24;
            end else begin
              roundCounter <= 4'h0;
            end
          end else begin
            if (_T_19) begin
              roundCounter <= 4'h0;
            end else begin
              if (io_en) begin
                roundCounter <= _T_24;
              end else begin
                roundCounter <= 4'h0;
              end
            end
          end
        end
      end else begin
        if (io_en) begin
          roundCounter <= _T_24;
        end else begin
          roundCounter <= 4'h0;
        end
      end
    end
    if (reset) begin
      state <= 128'h0;
    end else begin
      if (io_en) begin
        if (_T_396) begin
          state <= t;
        end else begin
          if (_T_401) begin
            state <= state3;
          end else begin
            state <= state31;
          end
        end
      end else begin
        state <= state31;
      end
    end
  end
endmodule
module expander( // @[:@1684.2]
  input          clock, // @[:@1685.4]
  input          reset, // @[:@1686.4]
  output [31:0]  io_sboxio_addr, // @[:@1687.4]
  input  [31:0]  io_sboxio_data, // @[:@1687.4]
  input  [3:0]   io_round, // @[:@1687.4]
  output [127:0] io_data, // @[:@1687.4]
  input  [127:0] io_key // @[:@1687.4]
);
  reg [127:0] pKey; // @[KeyExpander.scala 23:21:@1689.4]
  reg [127:0] _RAND_0;
  reg  gDone; // @[KeyExpander.scala 24:22:@1690.4]
  reg [31:0] _RAND_1;
  reg [127:0] roundkeys_0; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_2;
  reg [127:0] roundkeys_1; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_3;
  reg [127:0] roundkeys_2; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_4;
  reg [127:0] roundkeys_3; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_5;
  reg [127:0] roundkeys_4; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_6;
  reg [127:0] roundkeys_5; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_7;
  reg [127:0] roundkeys_6; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_8;
  reg [127:0] roundkeys_7; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_9;
  reg [127:0] roundkeys_8; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_10;
  reg [127:0] roundkeys_9; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_11;
  reg [127:0] roundkeys_10; // @[KeyExpander.scala 28:22:@1705.4]
  reg [127:0] _RAND_12;
  wire  _T_187; // @[KeyExpander.scala 117:22:@1770.6]
  wire [3:0] _GEN_93; // @[KeyExpander.scala 118:5:@1771.6]
  wire [3:0] tround; // @[KeyExpander.scala 93:5:@1758.4]
  wire [4:0] _T_143; // @[KeyExpander.scala 50:30:@1722.4]
  wire [4:0] _T_144; // @[KeyExpander.scala 50:30:@1723.4]
  wire [3:0] _T_145; // @[KeyExpander.scala 50:30:@1724.4]
  wire [127:0] _GEN_9; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_10; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_11; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_12; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_13; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_14; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_15; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_16; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_17; // @[KeyExpander.scala 51:20:@1725.4]
  wire [127:0] _GEN_18; // @[KeyExpander.scala 51:20:@1725.4]
  wire [31:0] prklast; // @[KeyExpander.scala 51:20:@1725.4]
  wire [23:0] _T_149; // @[KeyExpander.scala 53:24:@1726.4]
  wire [7:0] _T_150; // @[KeyExpander.scala 53:38:@1727.4]
  wire [31:0] rtw; // @[Cat.scala 30:58:@1728.4]
  wire [6:0] _GEN_121; // @[KeyExpander.scala 60:20:@1730.4]
  wire [6:0] rnd; // @[KeyExpander.scala 60:20:@1730.4]
  wire [4:0] _T_152; // @[KeyExpander.scala 61:28:@1731.4]
  wire [5:0] _T_154; // @[KeyExpander.scala 61:32:@1732.4]
  wire [5:0] _T_155; // @[KeyExpander.scala 61:32:@1733.4]
  wire [4:0] _T_156; // @[KeyExpander.scala 61:32:@1734.4]
  wire [3:0] _T_158; // @[:@1735.4]
  wire [7:0] _GEN_19; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_20; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_21; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_22; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_23; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_24; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_25; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_26; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_27; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_28; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_29; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_30; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_31; // @[Cat.scala 30:58:@1736.4]
  wire [7:0] _GEN_32; // @[Cat.scala 30:58:@1736.4]
  wire [31:0] rconw; // @[Cat.scala 30:58:@1736.4]
  wire [31:0] fk; // @[KeyExpander.scala 63:18:@1737.4]
  wire [31:0] _T_160; // @[KeyExpander.scala 66:20:@1738.4]
  wire [31:0] k0; // @[KeyExpander.scala 66:15:@1739.4]
  wire [31:0] _T_161; // @[KeyExpander.scala 67:20:@1740.4]
  wire [31:0] k1; // @[KeyExpander.scala 67:15:@1741.4]
  wire [31:0] _T_162; // @[KeyExpander.scala 68:20:@1742.4]
  wire [31:0] k2; // @[KeyExpander.scala 68:15:@1743.4]
  wire [31:0] k3; // @[KeyExpander.scala 69:15:@1745.4]
  wire [63:0] _T_164; // @[Cat.scala 30:58:@1746.4]
  wire [63:0] _T_165; // @[Cat.scala 30:58:@1747.4]
  wire [127:0] out; // @[Cat.scala 30:58:@1748.4]
  wire  _T_166; // @[KeyExpander.scala 75:18:@1749.4]
  wire [127:0] _GEN_33; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_34; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_35; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_36; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_37; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_38; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_39; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_40; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_41; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _GEN_42; // @[KeyExpander.scala 75:10:@1750.4]
  wire [127:0] _T_171; // @[KeyExpander.scala 75:10:@1750.4]
  wire  _T_173; // @[KeyExpander.scala 76:18:@1751.4]
  wire [127:0] _T_174; // @[KeyExpander.scala 76:10:@1752.4]
  wire [127:0] _T_175; // @[KeyExpander.scala 74:17:@1753.4]
  wire  _T_182; // @[Conditional.scala 37:30:@1760.6]
  wire  _GEN_43; // @[Conditional.scala 40:58:@1761.6]
  wire [127:0] _GEN_46; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_47; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_48; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_49; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_50; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_51; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_52; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_53; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_54; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_55; // @[KeyExpander.scala 133:29:@1786.10]
  wire [127:0] _GEN_56; // @[KeyExpander.scala 133:29:@1786.10]
  wire  _T_202; // @[KeyExpander.scala 136:25:@1790.10]
  wire [127:0] _GEN_57; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_58; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_59; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_60; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_61; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_62; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_63; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_64; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_65; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_66; // @[KeyExpander.scala 161:29:@1792.12]
  wire [127:0] _GEN_67; // @[KeyExpander.scala 161:29:@1792.12]
  wire  _T_207; // @[KeyExpander.scala 168:31:@1793.12]
  wire [127:0] _GEN_68; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_69; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_70; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_71; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_72; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_73; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_74; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_75; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_76; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_77; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_78; // @[KeyExpander.scala 136:31:@1791.10]
  wire  _GEN_79; // @[KeyExpander.scala 136:31:@1791.10]
  wire [127:0] _GEN_80; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_81; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_82; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_83; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_84; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_85; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_86; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_87; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_88; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_89; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_90; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_91; // @[KeyExpander.scala 132:7:@1785.8]
  wire  _GEN_92; // @[KeyExpander.scala 132:7:@1785.8]
  wire [127:0] _GEN_94; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_95; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_96; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_97; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_98; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_99; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_100; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_101; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_102; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_103; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_104; // @[KeyExpander.scala 118:5:@1771.6]
  wire [127:0] _GEN_105; // @[KeyExpander.scala 118:5:@1771.6]
  wire  _GEN_106; // @[KeyExpander.scala 118:5:@1771.6]
  wire  _GEN_107; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_109; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_110; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_111; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_112; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_113; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_114; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_115; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_116; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_117; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_118; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_119; // @[KeyExpander.scala 93:5:@1758.4]
  wire [127:0] _GEN_120; // @[KeyExpander.scala 93:5:@1758.4]
  assign _T_187 = gDone == 1'h0; // @[KeyExpander.scala 117:22:@1770.6]
  assign _GEN_93 = _T_187 ? io_round : 4'h0; // @[KeyExpander.scala 118:5:@1771.6]
  assign tround = gDone ? 4'h0 : _GEN_93; // @[KeyExpander.scala 93:5:@1758.4]
  assign _T_143 = tround - 4'h1; // @[KeyExpander.scala 50:30:@1722.4]
  assign _T_144 = $unsigned(_T_143); // @[KeyExpander.scala 50:30:@1723.4]
  assign _T_145 = _T_144[3:0]; // @[KeyExpander.scala 50:30:@1724.4]
  assign _GEN_9 = 4'h1 == _T_145 ? roundkeys_1 : roundkeys_0; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_10 = 4'h2 == _T_145 ? roundkeys_2 : _GEN_9; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_11 = 4'h3 == _T_145 ? roundkeys_3 : _GEN_10; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_12 = 4'h4 == _T_145 ? roundkeys_4 : _GEN_11; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_13 = 4'h5 == _T_145 ? roundkeys_5 : _GEN_12; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_14 = 4'h6 == _T_145 ? roundkeys_6 : _GEN_13; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_15 = 4'h7 == _T_145 ? roundkeys_7 : _GEN_14; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_16 = 4'h8 == _T_145 ? roundkeys_8 : _GEN_15; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_17 = 4'h9 == _T_145 ? roundkeys_9 : _GEN_16; // @[KeyExpander.scala 51:20:@1725.4]
  assign _GEN_18 = 4'ha == _T_145 ? roundkeys_10 : _GEN_17; // @[KeyExpander.scala 51:20:@1725.4]
  assign prklast = _GEN_18[31:0]; // @[KeyExpander.scala 51:20:@1725.4]
  assign _T_149 = prklast[23:0]; // @[KeyExpander.scala 53:24:@1726.4]
  assign _T_150 = prklast[31:24]; // @[KeyExpander.scala 53:38:@1727.4]
  assign rtw = {_T_149,_T_150}; // @[Cat.scala 30:58:@1728.4]
  assign _GEN_121 = {{3'd0}, tround}; // @[KeyExpander.scala 60:20:@1730.4]
  assign rnd = _GEN_121 << 2'h2; // @[KeyExpander.scala 60:20:@1730.4]
  assign _T_152 = rnd[6:2]; // @[KeyExpander.scala 61:28:@1731.4]
  assign _T_154 = _T_152 - 5'h1; // @[KeyExpander.scala 61:32:@1732.4]
  assign _T_155 = $unsigned(_T_154); // @[KeyExpander.scala 61:32:@1733.4]
  assign _T_156 = _T_155[4:0]; // @[KeyExpander.scala 61:32:@1734.4]
  assign _T_158 = _T_156[3:0]; // @[:@1735.4]
  assign _GEN_19 = 4'h1 == _T_158 ? 8'h2 : 8'h1; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_20 = 4'h2 == _T_158 ? 8'h4 : _GEN_19; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_21 = 4'h3 == _T_158 ? 8'h8 : _GEN_20; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_22 = 4'h4 == _T_158 ? 8'h10 : _GEN_21; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_23 = 4'h5 == _T_158 ? 8'h20 : _GEN_22; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_24 = 4'h6 == _T_158 ? 8'h40 : _GEN_23; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_25 = 4'h7 == _T_158 ? 8'h80 : _GEN_24; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_26 = 4'h8 == _T_158 ? 8'h1b : _GEN_25; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_27 = 4'h9 == _T_158 ? 8'h36 : _GEN_26; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_28 = 4'ha == _T_158 ? 8'h6c : _GEN_27; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_29 = 4'hb == _T_158 ? 8'hd8 : _GEN_28; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_30 = 4'hc == _T_158 ? 8'hab : _GEN_29; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_31 = 4'hd == _T_158 ? 8'h4d : _GEN_30; // @[Cat.scala 30:58:@1736.4]
  assign _GEN_32 = 4'he == _T_158 ? 8'h9a : _GEN_31; // @[Cat.scala 30:58:@1736.4]
  assign rconw = {_GEN_32,24'h0}; // @[Cat.scala 30:58:@1736.4]
  assign fk = rconw ^ io_sboxio_data; // @[KeyExpander.scala 63:18:@1737.4]
  assign _T_160 = _GEN_18[127:96]; // @[KeyExpander.scala 66:20:@1738.4]
  assign k0 = fk ^ _T_160; // @[KeyExpander.scala 66:15:@1739.4]
  assign _T_161 = _GEN_18[95:64]; // @[KeyExpander.scala 67:20:@1740.4]
  assign k1 = k0 ^ _T_161; // @[KeyExpander.scala 67:15:@1741.4]
  assign _T_162 = _GEN_18[63:32]; // @[KeyExpander.scala 68:20:@1742.4]
  assign k2 = k1 ^ _T_162; // @[KeyExpander.scala 68:15:@1743.4]
  assign k3 = k2 ^ prklast; // @[KeyExpander.scala 69:15:@1745.4]
  assign _T_164 = {k2,k3}; // @[Cat.scala 30:58:@1746.4]
  assign _T_165 = {k0,k1}; // @[Cat.scala 30:58:@1747.4]
  assign out = {_T_165,_T_164}; // @[Cat.scala 30:58:@1748.4]
  assign _T_166 = io_key == pKey; // @[KeyExpander.scala 75:18:@1749.4]
  assign _GEN_33 = 4'h1 == io_round ? roundkeys_1 : roundkeys_0; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_34 = 4'h2 == io_round ? roundkeys_2 : _GEN_33; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_35 = 4'h3 == io_round ? roundkeys_3 : _GEN_34; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_36 = 4'h4 == io_round ? roundkeys_4 : _GEN_35; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_37 = 4'h5 == io_round ? roundkeys_5 : _GEN_36; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_38 = 4'h6 == io_round ? roundkeys_6 : _GEN_37; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_39 = 4'h7 == io_round ? roundkeys_7 : _GEN_38; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_40 = 4'h8 == io_round ? roundkeys_8 : _GEN_39; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_41 = 4'h9 == io_round ? roundkeys_9 : _GEN_40; // @[KeyExpander.scala 75:10:@1750.4]
  assign _GEN_42 = 4'ha == io_round ? roundkeys_10 : _GEN_41; // @[KeyExpander.scala 75:10:@1750.4]
  assign _T_171 = _T_166 ? _GEN_42 : 128'h0; // @[KeyExpander.scala 75:10:@1750.4]
  assign _T_173 = tround == 4'h0; // @[KeyExpander.scala 76:18:@1751.4]
  assign _T_174 = _T_173 ? io_key : out; // @[KeyExpander.scala 76:10:@1752.4]
  assign _T_175 = gDone ? _T_171 : _T_174; // @[KeyExpander.scala 74:17:@1753.4]
  assign _T_182 = 1'h0 == _T_166; // @[Conditional.scala 37:30:@1760.6]
  assign _GEN_43 = _T_182 ? 1'h0 : gDone; // @[Conditional.scala 40:58:@1761.6]
  assign _GEN_46 = 4'h0 == tround ? io_key : roundkeys_0; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_47 = 4'h1 == tround ? io_key : roundkeys_1; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_48 = 4'h2 == tround ? io_key : roundkeys_2; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_49 = 4'h3 == tround ? io_key : roundkeys_3; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_50 = 4'h4 == tround ? io_key : roundkeys_4; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_51 = 4'h5 == tround ? io_key : roundkeys_5; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_52 = 4'h6 == tround ? io_key : roundkeys_6; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_53 = 4'h7 == tround ? io_key : roundkeys_7; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_54 = 4'h8 == tround ? io_key : roundkeys_8; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_55 = 4'h9 == tround ? io_key : roundkeys_9; // @[KeyExpander.scala 133:29:@1786.10]
  assign _GEN_56 = 4'ha == tround ? io_key : roundkeys_10; // @[KeyExpander.scala 133:29:@1786.10]
  assign _T_202 = tround > 4'h0; // @[KeyExpander.scala 136:25:@1790.10]
  assign _GEN_57 = 4'h0 == tround ? out : roundkeys_0; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_58 = 4'h1 == tround ? out : roundkeys_1; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_59 = 4'h2 == tround ? out : roundkeys_2; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_60 = 4'h3 == tround ? out : roundkeys_3; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_61 = 4'h4 == tround ? out : roundkeys_4; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_62 = 4'h5 == tround ? out : roundkeys_5; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_63 = 4'h6 == tround ? out : roundkeys_6; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_64 = 4'h7 == tround ? out : roundkeys_7; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_65 = 4'h8 == tround ? out : roundkeys_8; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_66 = 4'h9 == tround ? out : roundkeys_9; // @[KeyExpander.scala 161:29:@1792.12]
  assign _GEN_67 = 4'ha == tround ? out : roundkeys_10; // @[KeyExpander.scala 161:29:@1792.12]
  assign _T_207 = tround == 4'ha; // @[KeyExpander.scala 168:31:@1793.12]
  assign _GEN_68 = _T_202 ? _GEN_57 : roundkeys_0; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_69 = _T_202 ? _GEN_58 : roundkeys_1; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_70 = _T_202 ? _GEN_59 : roundkeys_2; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_71 = _T_202 ? _GEN_60 : roundkeys_3; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_72 = _T_202 ? _GEN_61 : roundkeys_4; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_73 = _T_202 ? _GEN_62 : roundkeys_5; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_74 = _T_202 ? _GEN_63 : roundkeys_6; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_75 = _T_202 ? _GEN_64 : roundkeys_7; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_76 = _T_202 ? _GEN_65 : roundkeys_8; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_77 = _T_202 ? _GEN_66 : roundkeys_9; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_78 = _T_202 ? _GEN_67 : roundkeys_10; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_79 = _T_202 ? _T_207 : gDone; // @[KeyExpander.scala 136:31:@1791.10]
  assign _GEN_80 = _T_173 ? _GEN_46 : _GEN_68; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_81 = _T_173 ? _GEN_47 : _GEN_69; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_82 = _T_173 ? _GEN_48 : _GEN_70; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_83 = _T_173 ? _GEN_49 : _GEN_71; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_84 = _T_173 ? _GEN_50 : _GEN_72; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_85 = _T_173 ? _GEN_51 : _GEN_73; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_86 = _T_173 ? _GEN_52 : _GEN_74; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_87 = _T_173 ? _GEN_53 : _GEN_75; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_88 = _T_173 ? _GEN_54 : _GEN_76; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_89 = _T_173 ? _GEN_55 : _GEN_77; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_90 = _T_173 ? _GEN_56 : _GEN_78; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_91 = _T_173 ? io_key : pKey; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_92 = _T_173 ? gDone : _GEN_79; // @[KeyExpander.scala 132:7:@1785.8]
  assign _GEN_94 = _T_187 ? _GEN_80 : roundkeys_0; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_95 = _T_187 ? _GEN_81 : roundkeys_1; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_96 = _T_187 ? _GEN_82 : roundkeys_2; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_97 = _T_187 ? _GEN_83 : roundkeys_3; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_98 = _T_187 ? _GEN_84 : roundkeys_4; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_99 = _T_187 ? _GEN_85 : roundkeys_5; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_100 = _T_187 ? _GEN_86 : roundkeys_6; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_101 = _T_187 ? _GEN_87 : roundkeys_7; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_102 = _T_187 ? _GEN_88 : roundkeys_8; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_103 = _T_187 ? _GEN_89 : roundkeys_9; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_104 = _T_187 ? _GEN_90 : roundkeys_10; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_105 = _T_187 ? _GEN_91 : pKey; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_106 = _T_187 ? _GEN_92 : gDone; // @[KeyExpander.scala 118:5:@1771.6]
  assign _GEN_107 = gDone ? _GEN_43 : _GEN_106; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_109 = gDone ? roundkeys_0 : _GEN_94; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_110 = gDone ? roundkeys_1 : _GEN_95; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_111 = gDone ? roundkeys_2 : _GEN_96; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_112 = gDone ? roundkeys_3 : _GEN_97; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_113 = gDone ? roundkeys_4 : _GEN_98; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_114 = gDone ? roundkeys_5 : _GEN_99; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_115 = gDone ? roundkeys_6 : _GEN_100; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_116 = gDone ? roundkeys_7 : _GEN_101; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_117 = gDone ? roundkeys_8 : _GEN_102; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_118 = gDone ? roundkeys_9 : _GEN_103; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_119 = gDone ? roundkeys_10 : _GEN_104; // @[KeyExpander.scala 93:5:@1758.4]
  assign _GEN_120 = gDone ? pKey : _GEN_105; // @[KeyExpander.scala 93:5:@1758.4]
  assign io_sboxio_addr = rtw;
  assign io_data = _T_175;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{$random}};
  pKey = _RAND_0[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  gDone = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {4{$random}};
  roundkeys_0 = _RAND_2[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {4{$random}};
  roundkeys_1 = _RAND_3[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {4{$random}};
  roundkeys_2 = _RAND_4[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {4{$random}};
  roundkeys_3 = _RAND_5[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {4{$random}};
  roundkeys_4 = _RAND_6[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {4{$random}};
  roundkeys_5 = _RAND_7[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {4{$random}};
  roundkeys_6 = _RAND_8[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {4{$random}};
  roundkeys_7 = _RAND_9[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {4{$random}};
  roundkeys_8 = _RAND_10[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {4{$random}};
  roundkeys_9 = _RAND_11[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {4{$random}};
  roundkeys_10 = _RAND_12[127:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pKey <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            pKey <= io_key;
          end
        end
      end
    end
    if (reset) begin
      gDone <= 1'h0;
    end else begin
      if (gDone) begin
        if (_T_182) begin
          gDone <= 1'h0;
        end
      end else begin
        if (_T_187) begin
          if (!(_T_173)) begin
            if (_T_202) begin
              gDone <= _T_207;
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_0 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h0 == tround) begin
              roundkeys_0 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h0 == tround) begin
                roundkeys_0 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_1 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h1 == tround) begin
              roundkeys_1 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h1 == tround) begin
                roundkeys_1 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_2 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h2 == tround) begin
              roundkeys_2 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h2 == tround) begin
                roundkeys_2 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_3 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h3 == tround) begin
              roundkeys_3 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h3 == tround) begin
                roundkeys_3 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_4 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h4 == tround) begin
              roundkeys_4 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h4 == tround) begin
                roundkeys_4 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_5 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h5 == tround) begin
              roundkeys_5 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h5 == tround) begin
                roundkeys_5 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_6 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h6 == tround) begin
              roundkeys_6 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h6 == tround) begin
                roundkeys_6 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_7 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h7 == tround) begin
              roundkeys_7 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h7 == tround) begin
                roundkeys_7 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_8 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h8 == tround) begin
              roundkeys_8 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h8 == tround) begin
                roundkeys_8 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_9 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'h9 == tround) begin
              roundkeys_9 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'h9 == tround) begin
                roundkeys_9 <= out;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      roundkeys_10 <= 128'h0;
    end else begin
      if (!(gDone)) begin
        if (_T_187) begin
          if (_T_173) begin
            if (4'ha == tround) begin
              roundkeys_10 <= io_key;
            end
          end else begin
            if (_T_202) begin
              if (4'ha == tround) begin
                roundkeys_10 <= out;
              end
            end
          end
        end
      end
    end
  end
endmodule
module sbox( // @[:@1799.2]
  input  [31:0]  io_addr, // @[:@1802.4]
  output [31:0]  io_data, // @[:@1802.4]
  input  [127:0] io_addr2, // @[:@1802.4]
  output [127:0] io_data2 // @[:@1802.4]
);
  wire [7:0] _T_522; // @[sbox.scala 46:24:@2061.4]
  wire [7:0] _T_524; // @[sbox.scala 47:24:@2062.4]
  wire [7:0] _T_526; // @[sbox.scala 48:24:@2063.4]
  wire [7:0] _T_528; // @[sbox.scala 49:24:@2064.4]
  wire [7:0] _GEN_20; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_21; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_22; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_23; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_24; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_25; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_26; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_27; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_28; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_29; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_30; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_31; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_32; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_33; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_34; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_35; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_36; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_37; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_38; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_39; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_40; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_41; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_42; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_43; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_44; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_45; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_46; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_47; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_48; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_49; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_50; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_51; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_52; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_53; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_54; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_55; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_56; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_57; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_58; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_59; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_60; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_61; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_62; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_63; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_64; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_65; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_66; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_67; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_68; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_69; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_70; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_71; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_72; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_73; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_74; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_75; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_76; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_77; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_78; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_79; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_80; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_81; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_82; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_83; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_84; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_85; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_86; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_87; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_88; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_89; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_90; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_91; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_92; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_93; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_94; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_95; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_96; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_97; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_98; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_99; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_100; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_101; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_102; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_103; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_104; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_105; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_106; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_107; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_108; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_109; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_110; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_111; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_112; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_113; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_114; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_115; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_116; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_117; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_118; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_119; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_120; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_121; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_122; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_123; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_124; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_125; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_126; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_127; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_128; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_129; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_130; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_131; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_132; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_133; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_134; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_135; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_136; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_137; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_138; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_139; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_140; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_141; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_142; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_143; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_144; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_145; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_146; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_147; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_148; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_149; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_150; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_151; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_152; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_153; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_154; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_155; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_156; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_157; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_158; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_159; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_160; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_161; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_162; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_163; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_164; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_165; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_166; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_167; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_168; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_169; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_170; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_171; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_172; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_173; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_174; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_175; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_176; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_177; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_178; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_179; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_180; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_181; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_182; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_183; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_184; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_185; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_186; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_187; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_188; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_189; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_190; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_191; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_192; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_193; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_194; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_195; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_196; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_197; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_198; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_199; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_200; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_201; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_202; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_203; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_204; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_205; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_206; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_207; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_208; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_209; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_210; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_211; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_212; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_213; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_214; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_215; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_216; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_217; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_218; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_219; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_220; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_221; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_222; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_223; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_224; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_225; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_226; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_227; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_228; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_229; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_230; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_231; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_232; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_233; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_234; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_235; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_236; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_237; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_238; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_239; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_240; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_241; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_242; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_243; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_244; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_245; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_246; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_247; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_248; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_249; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_250; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_251; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_252; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_253; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_254; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_255; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_256; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_257; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_258; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_259; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_260; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_261; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_262; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_263; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_264; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_265; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_266; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_267; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_268; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_269; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_270; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_271; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_272; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_273; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_274; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_275; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_276; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_277; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_278; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_279; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_280; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_281; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_282; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_283; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_284; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_285; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_286; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_287; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_288; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_289; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_290; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_291; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_292; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_293; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_294; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_295; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_296; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_297; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_298; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_299; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_300; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_301; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_302; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_303; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_304; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_305; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_306; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_307; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_308; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_309; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_310; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_311; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_312; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_313; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_314; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_315; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_316; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_317; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_318; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_319; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_320; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_321; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_322; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_323; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_324; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_325; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_326; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_327; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_328; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_329; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_330; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_331; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_332; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_333; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_334; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_335; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_336; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_337; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_338; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_339; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_340; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_341; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_342; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_343; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_344; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_345; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_346; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_347; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_348; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_349; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_350; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_351; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_352; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_353; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_354; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_355; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_356; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_357; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_358; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_359; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_360; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_361; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_362; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_363; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_364; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_365; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_366; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_367; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_368; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_369; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_370; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_371; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_372; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_373; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_374; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_375; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_376; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_377; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_378; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_379; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_380; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_381; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_382; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_383; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_384; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_385; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_386; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_387; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_388; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_389; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_390; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_391; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_392; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_393; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_394; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_395; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_396; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_397; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_398; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_399; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_400; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_401; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_402; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_403; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_404; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_405; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_406; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_407; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_408; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_409; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_410; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_411; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_412; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_413; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_414; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_415; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_416; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_417; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_418; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_419; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_420; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_421; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_422; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_423; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_424; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_425; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_426; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_427; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_428; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_429; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_430; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_431; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_432; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_433; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_434; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_435; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_436; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_437; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_438; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_439; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_440; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_441; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_442; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_443; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_444; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_445; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_446; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_447; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_448; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_449; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_450; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_451; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_452; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_453; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_454; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_455; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_456; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_457; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_458; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_459; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_460; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_461; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_462; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_463; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_464; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_465; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_466; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_467; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_468; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_469; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_470; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_471; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_472; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_473; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_474; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_475; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_476; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_477; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_478; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_479; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_480; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_481; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_482; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_483; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_484; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_485; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_486; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_487; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_488; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_489; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_490; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_491; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_492; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_493; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_494; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_495; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_496; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_497; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_498; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_499; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_500; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_501; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_502; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_503; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_504; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_505; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_506; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_507; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_508; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_509; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_510; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_511; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_512; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_513; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_514; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_515; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_516; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_517; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_518; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_519; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_520; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_521; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_522; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_523; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_524; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_525; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_526; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_527; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_528; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_529; // @[Cat.scala 30:58:@2065.4]
  wire [15:0] _T_530; // @[Cat.scala 30:58:@2065.4]
  wire [7:0] _GEN_530; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_531; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_532; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_533; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_534; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_535; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_536; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_537; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_538; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_539; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_540; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_541; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_542; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_543; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_544; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_545; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_546; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_547; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_548; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_549; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_550; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_551; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_552; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_553; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_554; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_555; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_556; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_557; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_558; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_559; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_560; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_561; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_562; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_563; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_564; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_565; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_566; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_567; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_568; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_569; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_570; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_571; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_572; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_573; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_574; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_575; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_576; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_577; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_578; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_579; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_580; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_581; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_582; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_583; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_584; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_585; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_586; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_587; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_588; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_589; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_590; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_591; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_592; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_593; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_594; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_595; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_596; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_597; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_598; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_599; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_600; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_601; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_602; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_603; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_604; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_605; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_606; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_607; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_608; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_609; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_610; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_611; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_612; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_613; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_614; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_615; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_616; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_617; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_618; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_619; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_620; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_621; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_622; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_623; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_624; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_625; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_626; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_627; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_628; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_629; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_630; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_631; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_632; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_633; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_634; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_635; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_636; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_637; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_638; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_639; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_640; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_641; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_642; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_643; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_644; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_645; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_646; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_647; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_648; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_649; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_650; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_651; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_652; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_653; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_654; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_655; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_656; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_657; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_658; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_659; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_660; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_661; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_662; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_663; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_664; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_665; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_666; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_667; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_668; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_669; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_670; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_671; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_672; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_673; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_674; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_675; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_676; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_677; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_678; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_679; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_680; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_681; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_682; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_683; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_684; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_685; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_686; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_687; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_688; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_689; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_690; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_691; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_692; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_693; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_694; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_695; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_696; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_697; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_698; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_699; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_700; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_701; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_702; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_703; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_704; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_705; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_706; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_707; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_708; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_709; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_710; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_711; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_712; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_713; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_714; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_715; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_716; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_717; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_718; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_719; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_720; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_721; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_722; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_723; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_724; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_725; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_726; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_727; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_728; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_729; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_730; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_731; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_732; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_733; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_734; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_735; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_736; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_737; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_738; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_739; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_740; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_741; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_742; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_743; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_744; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_745; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_746; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_747; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_748; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_749; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_750; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_751; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_752; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_753; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_754; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_755; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_756; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_757; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_758; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_759; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_760; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_761; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_762; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_763; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_764; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_765; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_766; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_767; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_768; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_769; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_770; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_771; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_772; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_773; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_774; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_775; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_776; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_777; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_778; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_779; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_780; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_781; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_782; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_783; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_784; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_785; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_786; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_787; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_788; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_789; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_790; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_791; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_792; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_793; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_794; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_795; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_796; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_797; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_798; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_799; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_800; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_801; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_802; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_803; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_804; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_805; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_806; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_807; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_808; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_809; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_810; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_811; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_812; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_813; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_814; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_815; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_816; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_817; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_818; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_819; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_820; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_821; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_822; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_823; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_824; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_825; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_826; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_827; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_828; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_829; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_830; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_831; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_832; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_833; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_834; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_835; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_836; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_837; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_838; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_839; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_840; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_841; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_842; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_843; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_844; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_845; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_846; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_847; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_848; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_849; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_850; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_851; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_852; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_853; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_854; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_855; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_856; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_857; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_858; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_859; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_860; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_861; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_862; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_863; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_864; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_865; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_866; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_867; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_868; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_869; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_870; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_871; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_872; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_873; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_874; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_875; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_876; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_877; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_878; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_879; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_880; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_881; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_882; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_883; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_884; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_885; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_886; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_887; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_888; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_889; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_890; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_891; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_892; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_893; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_894; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_895; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_896; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_897; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_898; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_899; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_900; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_901; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_902; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_903; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_904; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_905; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_906; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_907; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_908; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_909; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_910; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_911; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_912; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_913; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_914; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_915; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_916; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_917; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_918; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_919; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_920; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_921; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_922; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_923; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_924; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_925; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_926; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_927; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_928; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_929; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_930; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_931; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_932; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_933; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_934; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_935; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_936; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_937; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_938; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_939; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_940; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_941; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_942; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_943; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_944; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_945; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_946; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_947; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_948; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_949; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_950; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_951; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_952; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_953; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_954; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_955; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_956; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_957; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_958; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_959; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_960; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_961; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_962; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_963; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_964; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_965; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_966; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_967; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_968; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_969; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_970; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_971; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_972; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_973; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_974; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_975; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_976; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_977; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_978; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_979; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_980; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_981; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_982; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_983; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_984; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_985; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_986; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_987; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_988; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_989; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_990; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_991; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_992; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_993; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_994; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_995; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_996; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_997; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_998; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_999; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1000; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1001; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1002; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1003; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1004; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1005; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1006; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1007; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1008; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1009; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1010; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1011; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1012; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1013; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1014; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1015; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1016; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1017; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1018; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1019; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1020; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1021; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1022; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1023; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1024; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1025; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1026; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1027; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1028; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1029; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1030; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1031; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1032; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1033; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1034; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1035; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1036; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1037; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1038; // @[Cat.scala 30:58:@2066.4]
  wire [7:0] _GEN_1039; // @[Cat.scala 30:58:@2066.4]
  wire [15:0] _T_531; // @[Cat.scala 30:58:@2066.4]
  wire [31:0] _T_532; // @[Cat.scala 30:58:@2067.4]
  wire [7:0] _T_533; // @[sbox.scala 55:25:@2069.4]
  wire [7:0] _T_535; // @[sbox.scala 56:25:@2070.4]
  wire [7:0] _T_537; // @[sbox.scala 57:25:@2071.4]
  wire [7:0] _T_539; // @[sbox.scala 58:25:@2072.4]
  wire [7:0] _GEN_1040; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1041; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1042; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1043; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1044; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1045; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1046; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1047; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1048; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1049; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1050; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1051; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1052; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1053; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1054; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1055; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1056; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1057; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1058; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1059; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1060; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1061; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1062; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1063; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1064; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1065; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1066; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1067; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1068; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1069; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1070; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1071; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1072; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1073; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1074; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1075; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1076; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1077; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1078; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1079; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1080; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1081; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1082; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1083; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1084; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1085; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1086; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1087; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1088; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1089; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1090; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1091; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1092; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1093; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1094; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1095; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1096; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1097; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1098; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1099; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1100; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1101; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1102; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1103; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1104; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1105; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1106; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1107; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1108; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1109; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1110; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1111; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1112; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1113; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1114; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1115; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1116; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1117; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1118; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1119; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1120; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1121; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1122; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1123; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1124; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1125; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1126; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1127; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1128; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1129; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1130; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1131; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1132; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1133; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1134; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1135; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1136; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1137; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1138; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1139; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1140; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1141; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1142; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1143; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1144; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1145; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1146; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1147; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1148; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1149; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1150; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1151; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1152; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1153; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1154; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1155; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1156; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1157; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1158; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1159; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1160; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1161; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1162; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1163; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1164; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1165; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1166; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1167; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1168; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1169; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1170; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1171; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1172; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1173; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1174; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1175; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1176; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1177; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1178; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1179; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1180; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1181; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1182; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1183; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1184; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1185; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1186; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1187; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1188; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1189; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1190; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1191; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1192; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1193; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1194; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1195; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1196; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1197; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1198; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1199; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1200; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1201; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1202; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1203; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1204; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1205; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1206; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1207; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1208; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1209; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1210; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1211; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1212; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1213; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1214; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1215; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1216; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1217; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1218; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1219; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1220; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1221; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1222; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1223; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1224; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1225; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1226; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1227; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1228; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1229; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1230; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1231; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1232; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1233; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1234; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1235; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1236; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1237; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1238; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1239; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1240; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1241; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1242; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1243; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1244; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1245; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1246; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1247; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1248; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1249; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1250; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1251; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1252; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1253; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1254; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1255; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1256; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1257; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1258; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1259; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1260; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1261; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1262; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1263; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1264; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1265; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1266; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1267; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1268; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1269; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1270; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1271; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1272; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1273; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1274; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1275; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1276; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1277; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1278; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1279; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1280; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1281; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1282; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1283; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1284; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1285; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1286; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1287; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1288; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1289; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1290; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1291; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1292; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1293; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1294; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1295; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1296; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1297; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1298; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1299; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1300; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1301; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1302; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1303; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1304; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1305; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1306; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1307; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1308; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1309; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1310; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1311; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1312; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1313; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1314; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1315; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1316; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1317; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1318; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1319; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1320; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1321; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1322; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1323; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1324; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1325; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1326; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1327; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1328; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1329; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1330; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1331; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1332; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1333; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1334; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1335; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1336; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1337; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1338; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1339; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1340; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1341; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1342; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1343; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1344; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1345; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1346; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1347; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1348; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1349; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1350; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1351; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1352; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1353; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1354; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1355; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1356; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1357; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1358; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1359; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1360; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1361; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1362; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1363; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1364; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1365; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1366; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1367; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1368; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1369; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1370; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1371; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1372; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1373; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1374; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1375; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1376; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1377; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1378; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1379; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1380; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1381; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1382; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1383; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1384; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1385; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1386; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1387; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1388; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1389; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1390; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1391; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1392; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1393; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1394; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1395; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1396; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1397; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1398; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1399; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1400; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1401; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1402; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1403; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1404; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1405; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1406; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1407; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1408; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1409; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1410; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1411; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1412; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1413; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1414; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1415; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1416; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1417; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1418; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1419; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1420; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1421; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1422; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1423; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1424; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1425; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1426; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1427; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1428; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1429; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1430; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1431; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1432; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1433; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1434; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1435; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1436; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1437; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1438; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1439; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1440; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1441; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1442; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1443; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1444; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1445; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1446; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1447; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1448; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1449; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1450; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1451; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1452; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1453; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1454; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1455; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1456; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1457; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1458; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1459; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1460; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1461; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1462; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1463; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1464; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1465; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1466; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1467; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1468; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1469; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1470; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1471; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1472; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1473; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1474; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1475; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1476; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1477; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1478; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1479; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1480; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1481; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1482; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1483; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1484; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1485; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1486; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1487; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1488; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1489; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1490; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1491; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1492; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1493; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1494; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1495; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1496; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1497; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1498; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1499; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1500; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1501; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1502; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1503; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1504; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1505; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1506; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1507; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1508; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1509; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1510; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1511; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1512; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1513; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1514; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1515; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1516; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1517; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1518; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1519; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1520; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1521; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1522; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1523; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1524; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1525; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1526; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1527; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1528; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1529; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1530; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1531; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1532; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1533; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1534; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1535; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1536; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1537; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1538; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1539; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1540; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1541; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1542; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1543; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1544; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1545; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1546; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1547; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1548; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1549; // @[Cat.scala 30:58:@2073.4]
  wire [15:0] _T_541; // @[Cat.scala 30:58:@2073.4]
  wire [7:0] _GEN_1550; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1551; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1552; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1553; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1554; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1555; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1556; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1557; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1558; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1559; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1560; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1561; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1562; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1563; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1564; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1565; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1566; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1567; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1568; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1569; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1570; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1571; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1572; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1573; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1574; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1575; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1576; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1577; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1578; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1579; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1580; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1581; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1582; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1583; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1584; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1585; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1586; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1587; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1588; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1589; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1590; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1591; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1592; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1593; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1594; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1595; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1596; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1597; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1598; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1599; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1600; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1601; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1602; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1603; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1604; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1605; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1606; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1607; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1608; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1609; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1610; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1611; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1612; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1613; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1614; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1615; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1616; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1617; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1618; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1619; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1620; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1621; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1622; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1623; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1624; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1625; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1626; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1627; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1628; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1629; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1630; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1631; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1632; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1633; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1634; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1635; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1636; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1637; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1638; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1639; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1640; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1641; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1642; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1643; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1644; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1645; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1646; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1647; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1648; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1649; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1650; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1651; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1652; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1653; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1654; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1655; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1656; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1657; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1658; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1659; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1660; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1661; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1662; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1663; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1664; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1665; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1666; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1667; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1668; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1669; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1670; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1671; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1672; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1673; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1674; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1675; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1676; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1677; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1678; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1679; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1680; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1681; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1682; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1683; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1684; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1685; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1686; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1687; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1688; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1689; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1690; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1691; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1692; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1693; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1694; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1695; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1696; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1697; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1698; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1699; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1700; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1701; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1702; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1703; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1704; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1705; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1706; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1707; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1708; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1709; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1710; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1711; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1712; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1713; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1714; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1715; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1716; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1717; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1718; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1719; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1720; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1721; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1722; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1723; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1724; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1725; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1726; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1727; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1728; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1729; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1730; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1731; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1732; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1733; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1734; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1735; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1736; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1737; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1738; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1739; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1740; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1741; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1742; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1743; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1744; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1745; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1746; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1747; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1748; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1749; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1750; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1751; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1752; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1753; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1754; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1755; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1756; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1757; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1758; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1759; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1760; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1761; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1762; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1763; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1764; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1765; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1766; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1767; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1768; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1769; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1770; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1771; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1772; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1773; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1774; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1775; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1776; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1777; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1778; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1779; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1780; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1781; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1782; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1783; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1784; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1785; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1786; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1787; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1788; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1789; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1790; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1791; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1792; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1793; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1794; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1795; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1796; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1797; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1798; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1799; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1800; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1801; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1802; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1803; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1804; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1805; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1806; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1807; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1808; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1809; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1810; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1811; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1812; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1813; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1814; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1815; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1816; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1817; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1818; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1819; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1820; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1821; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1822; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1823; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1824; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1825; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1826; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1827; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1828; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1829; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1830; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1831; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1832; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1833; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1834; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1835; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1836; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1837; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1838; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1839; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1840; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1841; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1842; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1843; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1844; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1845; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1846; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1847; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1848; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1849; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1850; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1851; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1852; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1853; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1854; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1855; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1856; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1857; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1858; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1859; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1860; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1861; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1862; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1863; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1864; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1865; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1866; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1867; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1868; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1869; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1870; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1871; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1872; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1873; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1874; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1875; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1876; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1877; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1878; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1879; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1880; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1881; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1882; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1883; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1884; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1885; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1886; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1887; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1888; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1889; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1890; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1891; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1892; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1893; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1894; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1895; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1896; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1897; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1898; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1899; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1900; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1901; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1902; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1903; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1904; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1905; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1906; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1907; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1908; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1909; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1910; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1911; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1912; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1913; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1914; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1915; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1916; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1917; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1918; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1919; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1920; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1921; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1922; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1923; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1924; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1925; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1926; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1927; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1928; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1929; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1930; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1931; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1932; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1933; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1934; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1935; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1936; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1937; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1938; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1939; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1940; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1941; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1942; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1943; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1944; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1945; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1946; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1947; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1948; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1949; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1950; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1951; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1952; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1953; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1954; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1955; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1956; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1957; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1958; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1959; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1960; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1961; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1962; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1963; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1964; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1965; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1966; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1967; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1968; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1969; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1970; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1971; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1972; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1973; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1974; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1975; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1976; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1977; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1978; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1979; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1980; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1981; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1982; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1983; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1984; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1985; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1986; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1987; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1988; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1989; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1990; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1991; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1992; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1993; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1994; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1995; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1996; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1997; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1998; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_1999; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2000; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2001; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2002; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2003; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2004; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2005; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2006; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2007; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2008; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2009; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2010; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2011; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2012; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2013; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2014; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2015; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2016; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2017; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2018; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2019; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2020; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2021; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2022; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2023; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2024; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2025; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2026; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2027; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2028; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2029; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2030; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2031; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2032; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2033; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2034; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2035; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2036; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2037; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2038; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2039; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2040; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2041; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2042; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2043; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2044; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2045; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2046; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2047; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2048; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2049; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2050; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2051; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2052; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2053; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2054; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2055; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2056; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2057; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2058; // @[Cat.scala 30:58:@2074.4]
  wire [7:0] _GEN_2059; // @[Cat.scala 30:58:@2074.4]
  wire [15:0] _T_542; // @[Cat.scala 30:58:@2074.4]
  wire [31:0] x1; // @[Cat.scala 30:58:@2075.4]
  wire [7:0] _T_543; // @[sbox.scala 62:25:@2076.4]
  wire [7:0] _T_545; // @[sbox.scala 63:25:@2077.4]
  wire [7:0] _T_547; // @[sbox.scala 64:26:@2078.4]
  wire [7:0] _T_549; // @[sbox.scala 65:26:@2079.4]
  wire [7:0] _GEN_2060; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2061; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2062; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2063; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2064; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2065; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2066; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2067; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2068; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2069; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2070; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2071; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2072; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2073; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2074; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2075; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2076; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2077; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2078; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2079; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2080; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2081; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2082; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2083; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2084; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2085; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2086; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2087; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2088; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2089; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2090; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2091; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2092; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2093; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2094; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2095; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2096; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2097; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2098; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2099; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2100; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2101; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2102; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2103; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2104; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2105; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2106; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2107; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2108; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2109; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2110; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2111; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2112; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2113; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2114; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2115; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2116; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2117; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2118; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2119; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2120; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2121; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2122; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2123; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2124; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2125; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2126; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2127; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2128; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2129; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2130; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2131; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2132; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2133; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2134; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2135; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2136; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2137; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2138; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2139; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2140; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2141; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2142; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2143; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2144; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2145; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2146; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2147; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2148; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2149; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2150; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2151; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2152; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2153; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2154; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2155; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2156; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2157; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2158; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2159; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2160; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2161; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2162; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2163; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2164; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2165; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2166; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2167; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2168; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2169; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2170; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2171; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2172; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2173; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2174; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2175; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2176; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2177; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2178; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2179; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2180; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2181; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2182; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2183; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2184; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2185; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2186; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2187; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2188; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2189; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2190; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2191; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2192; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2193; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2194; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2195; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2196; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2197; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2198; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2199; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2200; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2201; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2202; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2203; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2204; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2205; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2206; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2207; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2208; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2209; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2210; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2211; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2212; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2213; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2214; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2215; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2216; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2217; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2218; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2219; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2220; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2221; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2222; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2223; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2224; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2225; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2226; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2227; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2228; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2229; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2230; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2231; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2232; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2233; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2234; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2235; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2236; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2237; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2238; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2239; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2240; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2241; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2242; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2243; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2244; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2245; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2246; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2247; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2248; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2249; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2250; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2251; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2252; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2253; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2254; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2255; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2256; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2257; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2258; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2259; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2260; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2261; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2262; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2263; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2264; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2265; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2266; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2267; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2268; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2269; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2270; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2271; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2272; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2273; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2274; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2275; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2276; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2277; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2278; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2279; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2280; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2281; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2282; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2283; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2284; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2285; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2286; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2287; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2288; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2289; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2290; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2291; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2292; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2293; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2294; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2295; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2296; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2297; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2298; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2299; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2300; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2301; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2302; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2303; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2304; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2305; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2306; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2307; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2308; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2309; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2310; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2311; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2312; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2313; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2314; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2315; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2316; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2317; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2318; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2319; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2320; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2321; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2322; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2323; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2324; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2325; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2326; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2327; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2328; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2329; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2330; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2331; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2332; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2333; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2334; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2335; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2336; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2337; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2338; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2339; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2340; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2341; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2342; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2343; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2344; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2345; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2346; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2347; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2348; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2349; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2350; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2351; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2352; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2353; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2354; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2355; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2356; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2357; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2358; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2359; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2360; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2361; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2362; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2363; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2364; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2365; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2366; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2367; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2368; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2369; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2370; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2371; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2372; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2373; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2374; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2375; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2376; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2377; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2378; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2379; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2380; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2381; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2382; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2383; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2384; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2385; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2386; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2387; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2388; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2389; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2390; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2391; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2392; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2393; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2394; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2395; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2396; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2397; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2398; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2399; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2400; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2401; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2402; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2403; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2404; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2405; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2406; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2407; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2408; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2409; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2410; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2411; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2412; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2413; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2414; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2415; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2416; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2417; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2418; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2419; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2420; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2421; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2422; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2423; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2424; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2425; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2426; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2427; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2428; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2429; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2430; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2431; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2432; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2433; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2434; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2435; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2436; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2437; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2438; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2439; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2440; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2441; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2442; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2443; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2444; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2445; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2446; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2447; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2448; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2449; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2450; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2451; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2452; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2453; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2454; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2455; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2456; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2457; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2458; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2459; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2460; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2461; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2462; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2463; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2464; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2465; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2466; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2467; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2468; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2469; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2470; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2471; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2472; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2473; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2474; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2475; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2476; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2477; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2478; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2479; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2480; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2481; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2482; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2483; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2484; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2485; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2486; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2487; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2488; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2489; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2490; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2491; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2492; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2493; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2494; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2495; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2496; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2497; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2498; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2499; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2500; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2501; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2502; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2503; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2504; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2505; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2506; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2507; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2508; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2509; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2510; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2511; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2512; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2513; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2514; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2515; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2516; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2517; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2518; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2519; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2520; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2521; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2522; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2523; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2524; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2525; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2526; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2527; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2528; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2529; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2530; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2531; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2532; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2533; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2534; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2535; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2536; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2537; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2538; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2539; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2540; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2541; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2542; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2543; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2544; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2545; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2546; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2547; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2548; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2549; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2550; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2551; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2552; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2553; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2554; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2555; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2556; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2557; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2558; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2559; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2560; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2561; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2562; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2563; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2564; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2565; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2566; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2567; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2568; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2569; // @[Cat.scala 30:58:@2080.4]
  wire [15:0] _T_551; // @[Cat.scala 30:58:@2080.4]
  wire [7:0] _GEN_2570; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2571; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2572; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2573; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2574; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2575; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2576; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2577; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2578; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2579; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2580; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2581; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2582; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2583; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2584; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2585; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2586; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2587; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2588; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2589; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2590; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2591; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2592; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2593; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2594; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2595; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2596; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2597; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2598; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2599; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2600; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2601; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2602; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2603; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2604; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2605; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2606; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2607; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2608; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2609; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2610; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2611; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2612; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2613; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2614; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2615; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2616; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2617; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2618; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2619; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2620; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2621; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2622; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2623; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2624; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2625; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2626; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2627; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2628; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2629; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2630; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2631; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2632; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2633; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2634; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2635; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2636; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2637; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2638; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2639; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2640; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2641; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2642; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2643; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2644; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2645; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2646; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2647; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2648; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2649; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2650; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2651; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2652; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2653; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2654; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2655; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2656; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2657; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2658; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2659; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2660; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2661; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2662; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2663; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2664; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2665; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2666; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2667; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2668; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2669; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2670; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2671; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2672; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2673; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2674; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2675; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2676; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2677; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2678; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2679; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2680; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2681; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2682; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2683; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2684; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2685; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2686; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2687; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2688; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2689; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2690; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2691; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2692; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2693; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2694; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2695; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2696; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2697; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2698; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2699; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2700; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2701; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2702; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2703; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2704; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2705; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2706; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2707; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2708; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2709; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2710; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2711; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2712; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2713; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2714; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2715; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2716; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2717; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2718; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2719; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2720; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2721; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2722; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2723; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2724; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2725; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2726; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2727; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2728; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2729; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2730; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2731; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2732; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2733; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2734; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2735; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2736; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2737; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2738; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2739; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2740; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2741; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2742; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2743; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2744; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2745; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2746; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2747; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2748; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2749; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2750; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2751; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2752; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2753; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2754; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2755; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2756; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2757; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2758; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2759; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2760; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2761; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2762; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2763; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2764; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2765; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2766; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2767; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2768; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2769; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2770; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2771; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2772; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2773; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2774; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2775; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2776; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2777; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2778; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2779; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2780; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2781; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2782; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2783; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2784; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2785; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2786; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2787; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2788; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2789; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2790; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2791; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2792; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2793; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2794; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2795; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2796; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2797; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2798; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2799; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2800; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2801; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2802; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2803; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2804; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2805; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2806; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2807; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2808; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2809; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2810; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2811; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2812; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2813; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2814; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2815; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2816; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2817; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2818; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2819; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2820; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2821; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2822; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2823; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2824; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2825; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2826; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2827; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2828; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2829; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2830; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2831; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2832; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2833; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2834; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2835; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2836; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2837; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2838; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2839; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2840; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2841; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2842; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2843; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2844; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2845; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2846; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2847; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2848; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2849; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2850; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2851; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2852; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2853; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2854; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2855; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2856; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2857; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2858; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2859; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2860; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2861; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2862; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2863; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2864; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2865; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2866; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2867; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2868; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2869; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2870; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2871; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2872; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2873; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2874; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2875; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2876; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2877; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2878; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2879; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2880; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2881; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2882; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2883; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2884; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2885; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2886; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2887; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2888; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2889; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2890; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2891; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2892; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2893; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2894; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2895; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2896; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2897; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2898; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2899; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2900; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2901; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2902; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2903; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2904; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2905; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2906; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2907; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2908; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2909; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2910; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2911; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2912; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2913; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2914; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2915; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2916; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2917; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2918; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2919; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2920; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2921; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2922; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2923; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2924; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2925; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2926; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2927; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2928; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2929; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2930; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2931; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2932; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2933; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2934; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2935; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2936; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2937; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2938; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2939; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2940; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2941; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2942; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2943; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2944; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2945; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2946; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2947; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2948; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2949; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2950; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2951; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2952; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2953; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2954; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2955; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2956; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2957; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2958; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2959; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2960; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2961; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2962; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2963; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2964; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2965; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2966; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2967; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2968; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2969; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2970; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2971; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2972; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2973; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2974; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2975; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2976; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2977; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2978; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2979; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2980; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2981; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2982; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2983; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2984; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2985; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2986; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2987; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2988; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2989; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2990; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2991; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2992; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2993; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2994; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2995; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2996; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2997; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2998; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_2999; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3000; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3001; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3002; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3003; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3004; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3005; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3006; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3007; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3008; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3009; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3010; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3011; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3012; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3013; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3014; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3015; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3016; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3017; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3018; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3019; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3020; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3021; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3022; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3023; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3024; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3025; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3026; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3027; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3028; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3029; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3030; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3031; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3032; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3033; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3034; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3035; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3036; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3037; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3038; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3039; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3040; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3041; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3042; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3043; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3044; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3045; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3046; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3047; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3048; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3049; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3050; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3051; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3052; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3053; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3054; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3055; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3056; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3057; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3058; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3059; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3060; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3061; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3062; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3063; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3064; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3065; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3066; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3067; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3068; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3069; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3070; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3071; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3072; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3073; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3074; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3075; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3076; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3077; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3078; // @[Cat.scala 30:58:@2081.4]
  wire [7:0] _GEN_3079; // @[Cat.scala 30:58:@2081.4]
  wire [15:0] _T_552; // @[Cat.scala 30:58:@2081.4]
  wire [31:0] x2; // @[Cat.scala 30:58:@2082.4]
  wire [7:0] _T_553; // @[sbox.scala 69:26:@2083.4]
  wire [7:0] _T_555; // @[sbox.scala 70:26:@2084.4]
  wire [7:0] _T_557; // @[sbox.scala 71:26:@2085.4]
  wire [7:0] _T_559; // @[sbox.scala 72:26:@2086.4]
  wire [7:0] _GEN_3080; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3081; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3082; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3083; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3084; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3085; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3086; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3087; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3088; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3089; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3090; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3091; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3092; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3093; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3094; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3095; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3096; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3097; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3098; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3099; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3100; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3101; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3102; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3103; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3104; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3105; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3106; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3107; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3108; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3109; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3110; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3111; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3112; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3113; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3114; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3115; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3116; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3117; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3118; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3119; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3120; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3121; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3122; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3123; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3124; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3125; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3126; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3127; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3128; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3129; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3130; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3131; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3132; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3133; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3134; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3135; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3136; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3137; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3138; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3139; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3140; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3141; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3142; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3143; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3144; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3145; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3146; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3147; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3148; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3149; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3150; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3151; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3152; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3153; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3154; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3155; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3156; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3157; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3158; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3159; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3160; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3161; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3162; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3163; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3164; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3165; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3166; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3167; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3168; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3169; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3170; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3171; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3172; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3173; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3174; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3175; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3176; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3177; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3178; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3179; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3180; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3181; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3182; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3183; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3184; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3185; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3186; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3187; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3188; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3189; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3190; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3191; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3192; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3193; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3194; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3195; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3196; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3197; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3198; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3199; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3200; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3201; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3202; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3203; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3204; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3205; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3206; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3207; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3208; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3209; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3210; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3211; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3212; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3213; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3214; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3215; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3216; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3217; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3218; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3219; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3220; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3221; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3222; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3223; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3224; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3225; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3226; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3227; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3228; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3229; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3230; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3231; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3232; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3233; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3234; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3235; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3236; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3237; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3238; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3239; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3240; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3241; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3242; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3243; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3244; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3245; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3246; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3247; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3248; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3249; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3250; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3251; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3252; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3253; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3254; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3255; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3256; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3257; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3258; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3259; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3260; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3261; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3262; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3263; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3264; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3265; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3266; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3267; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3268; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3269; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3270; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3271; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3272; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3273; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3274; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3275; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3276; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3277; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3278; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3279; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3280; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3281; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3282; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3283; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3284; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3285; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3286; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3287; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3288; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3289; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3290; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3291; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3292; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3293; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3294; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3295; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3296; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3297; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3298; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3299; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3300; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3301; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3302; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3303; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3304; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3305; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3306; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3307; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3308; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3309; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3310; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3311; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3312; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3313; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3314; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3315; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3316; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3317; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3318; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3319; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3320; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3321; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3322; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3323; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3324; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3325; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3326; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3327; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3328; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3329; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3330; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3331; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3332; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3333; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3334; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3335; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3336; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3337; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3338; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3339; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3340; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3341; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3342; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3343; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3344; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3345; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3346; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3347; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3348; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3349; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3350; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3351; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3352; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3353; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3354; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3355; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3356; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3357; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3358; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3359; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3360; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3361; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3362; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3363; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3364; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3365; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3366; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3367; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3368; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3369; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3370; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3371; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3372; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3373; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3374; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3375; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3376; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3377; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3378; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3379; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3380; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3381; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3382; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3383; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3384; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3385; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3386; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3387; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3388; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3389; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3390; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3391; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3392; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3393; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3394; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3395; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3396; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3397; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3398; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3399; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3400; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3401; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3402; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3403; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3404; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3405; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3406; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3407; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3408; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3409; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3410; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3411; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3412; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3413; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3414; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3415; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3416; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3417; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3418; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3419; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3420; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3421; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3422; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3423; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3424; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3425; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3426; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3427; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3428; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3429; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3430; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3431; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3432; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3433; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3434; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3435; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3436; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3437; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3438; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3439; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3440; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3441; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3442; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3443; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3444; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3445; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3446; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3447; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3448; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3449; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3450; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3451; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3452; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3453; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3454; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3455; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3456; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3457; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3458; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3459; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3460; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3461; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3462; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3463; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3464; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3465; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3466; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3467; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3468; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3469; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3470; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3471; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3472; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3473; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3474; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3475; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3476; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3477; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3478; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3479; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3480; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3481; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3482; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3483; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3484; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3485; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3486; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3487; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3488; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3489; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3490; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3491; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3492; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3493; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3494; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3495; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3496; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3497; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3498; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3499; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3500; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3501; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3502; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3503; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3504; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3505; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3506; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3507; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3508; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3509; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3510; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3511; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3512; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3513; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3514; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3515; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3516; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3517; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3518; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3519; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3520; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3521; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3522; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3523; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3524; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3525; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3526; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3527; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3528; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3529; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3530; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3531; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3532; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3533; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3534; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3535; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3536; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3537; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3538; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3539; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3540; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3541; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3542; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3543; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3544; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3545; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3546; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3547; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3548; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3549; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3550; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3551; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3552; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3553; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3554; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3555; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3556; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3557; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3558; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3559; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3560; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3561; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3562; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3563; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3564; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3565; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3566; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3567; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3568; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3569; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3570; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3571; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3572; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3573; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3574; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3575; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3576; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3577; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3578; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3579; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3580; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3581; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3582; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3583; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3584; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3585; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3586; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3587; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3588; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3589; // @[Cat.scala 30:58:@2087.4]
  wire [15:0] _T_561; // @[Cat.scala 30:58:@2087.4]
  wire [7:0] _GEN_3590; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3591; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3592; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3593; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3594; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3595; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3596; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3597; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3598; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3599; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3600; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3601; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3602; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3603; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3604; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3605; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3606; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3607; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3608; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3609; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3610; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3611; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3612; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3613; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3614; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3615; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3616; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3617; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3618; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3619; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3620; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3621; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3622; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3623; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3624; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3625; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3626; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3627; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3628; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3629; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3630; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3631; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3632; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3633; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3634; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3635; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3636; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3637; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3638; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3639; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3640; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3641; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3642; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3643; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3644; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3645; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3646; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3647; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3648; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3649; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3650; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3651; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3652; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3653; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3654; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3655; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3656; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3657; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3658; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3659; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3660; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3661; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3662; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3663; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3664; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3665; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3666; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3667; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3668; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3669; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3670; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3671; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3672; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3673; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3674; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3675; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3676; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3677; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3678; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3679; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3680; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3681; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3682; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3683; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3684; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3685; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3686; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3687; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3688; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3689; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3690; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3691; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3692; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3693; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3694; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3695; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3696; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3697; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3698; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3699; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3700; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3701; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3702; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3703; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3704; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3705; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3706; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3707; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3708; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3709; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3710; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3711; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3712; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3713; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3714; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3715; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3716; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3717; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3718; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3719; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3720; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3721; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3722; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3723; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3724; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3725; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3726; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3727; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3728; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3729; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3730; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3731; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3732; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3733; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3734; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3735; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3736; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3737; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3738; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3739; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3740; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3741; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3742; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3743; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3744; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3745; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3746; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3747; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3748; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3749; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3750; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3751; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3752; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3753; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3754; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3755; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3756; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3757; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3758; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3759; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3760; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3761; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3762; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3763; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3764; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3765; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3766; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3767; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3768; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3769; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3770; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3771; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3772; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3773; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3774; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3775; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3776; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3777; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3778; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3779; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3780; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3781; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3782; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3783; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3784; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3785; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3786; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3787; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3788; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3789; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3790; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3791; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3792; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3793; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3794; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3795; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3796; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3797; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3798; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3799; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3800; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3801; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3802; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3803; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3804; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3805; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3806; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3807; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3808; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3809; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3810; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3811; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3812; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3813; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3814; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3815; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3816; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3817; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3818; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3819; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3820; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3821; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3822; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3823; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3824; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3825; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3826; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3827; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3828; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3829; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3830; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3831; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3832; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3833; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3834; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3835; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3836; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3837; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3838; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3839; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3840; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3841; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3842; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3843; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3844; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3845; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3846; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3847; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3848; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3849; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3850; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3851; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3852; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3853; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3854; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3855; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3856; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3857; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3858; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3859; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3860; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3861; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3862; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3863; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3864; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3865; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3866; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3867; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3868; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3869; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3870; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3871; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3872; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3873; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3874; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3875; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3876; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3877; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3878; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3879; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3880; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3881; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3882; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3883; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3884; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3885; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3886; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3887; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3888; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3889; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3890; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3891; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3892; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3893; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3894; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3895; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3896; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3897; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3898; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3899; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3900; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3901; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3902; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3903; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3904; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3905; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3906; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3907; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3908; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3909; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3910; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3911; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3912; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3913; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3914; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3915; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3916; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3917; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3918; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3919; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3920; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3921; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3922; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3923; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3924; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3925; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3926; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3927; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3928; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3929; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3930; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3931; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3932; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3933; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3934; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3935; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3936; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3937; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3938; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3939; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3940; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3941; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3942; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3943; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3944; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3945; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3946; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3947; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3948; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3949; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3950; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3951; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3952; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3953; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3954; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3955; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3956; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3957; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3958; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3959; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3960; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3961; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3962; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3963; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3964; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3965; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3966; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3967; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3968; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3969; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3970; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3971; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3972; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3973; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3974; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3975; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3976; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3977; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3978; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3979; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3980; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3981; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3982; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3983; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3984; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3985; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3986; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3987; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3988; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3989; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3990; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3991; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3992; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3993; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3994; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3995; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3996; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3997; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3998; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_3999; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4000; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4001; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4002; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4003; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4004; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4005; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4006; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4007; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4008; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4009; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4010; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4011; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4012; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4013; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4014; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4015; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4016; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4017; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4018; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4019; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4020; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4021; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4022; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4023; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4024; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4025; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4026; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4027; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4028; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4029; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4030; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4031; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4032; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4033; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4034; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4035; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4036; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4037; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4038; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4039; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4040; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4041; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4042; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4043; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4044; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4045; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4046; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4047; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4048; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4049; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4050; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4051; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4052; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4053; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4054; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4055; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4056; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4057; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4058; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4059; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4060; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4061; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4062; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4063; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4064; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4065; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4066; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4067; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4068; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4069; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4070; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4071; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4072; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4073; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4074; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4075; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4076; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4077; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4078; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4079; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4080; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4081; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4082; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4083; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4084; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4085; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4086; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4087; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4088; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4089; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4090; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4091; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4092; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4093; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4094; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4095; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4096; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4097; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4098; // @[Cat.scala 30:58:@2088.4]
  wire [7:0] _GEN_4099; // @[Cat.scala 30:58:@2088.4]
  wire [15:0] _T_562; // @[Cat.scala 30:58:@2088.4]
  wire [31:0] x3; // @[Cat.scala 30:58:@2089.4]
  wire [7:0] _T_563; // @[sbox.scala 76:26:@2090.4]
  wire [7:0] _T_565; // @[sbox.scala 77:26:@2091.4]
  wire [7:0] _T_567; // @[sbox.scala 78:26:@2092.4]
  wire [7:0] _T_569; // @[sbox.scala 79:26:@2093.4]
  wire [7:0] _GEN_4100; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4101; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4102; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4103; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4104; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4105; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4106; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4107; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4108; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4109; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4110; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4111; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4112; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4113; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4114; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4115; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4116; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4117; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4118; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4119; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4120; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4121; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4122; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4123; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4124; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4125; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4126; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4127; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4128; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4129; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4130; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4131; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4132; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4133; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4134; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4135; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4136; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4137; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4138; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4139; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4140; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4141; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4142; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4143; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4144; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4145; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4146; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4147; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4148; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4149; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4150; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4151; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4152; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4153; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4154; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4155; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4156; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4157; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4158; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4159; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4160; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4161; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4162; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4163; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4164; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4165; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4166; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4167; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4168; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4169; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4170; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4171; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4172; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4173; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4174; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4175; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4176; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4177; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4178; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4179; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4180; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4181; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4182; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4183; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4184; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4185; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4186; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4187; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4188; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4189; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4190; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4191; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4192; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4193; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4194; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4195; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4196; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4197; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4198; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4199; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4200; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4201; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4202; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4203; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4204; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4205; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4206; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4207; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4208; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4209; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4210; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4211; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4212; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4213; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4214; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4215; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4216; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4217; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4218; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4219; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4220; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4221; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4222; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4223; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4224; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4225; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4226; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4227; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4228; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4229; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4230; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4231; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4232; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4233; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4234; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4235; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4236; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4237; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4238; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4239; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4240; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4241; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4242; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4243; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4244; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4245; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4246; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4247; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4248; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4249; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4250; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4251; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4252; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4253; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4254; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4255; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4256; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4257; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4258; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4259; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4260; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4261; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4262; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4263; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4264; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4265; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4266; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4267; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4268; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4269; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4270; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4271; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4272; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4273; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4274; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4275; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4276; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4277; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4278; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4279; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4280; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4281; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4282; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4283; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4284; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4285; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4286; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4287; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4288; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4289; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4290; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4291; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4292; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4293; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4294; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4295; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4296; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4297; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4298; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4299; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4300; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4301; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4302; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4303; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4304; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4305; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4306; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4307; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4308; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4309; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4310; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4311; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4312; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4313; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4314; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4315; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4316; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4317; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4318; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4319; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4320; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4321; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4322; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4323; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4324; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4325; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4326; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4327; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4328; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4329; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4330; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4331; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4332; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4333; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4334; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4335; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4336; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4337; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4338; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4339; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4340; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4341; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4342; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4343; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4344; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4345; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4346; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4347; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4348; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4349; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4350; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4351; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4352; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4353; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4354; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4355; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4356; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4357; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4358; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4359; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4360; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4361; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4362; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4363; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4364; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4365; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4366; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4367; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4368; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4369; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4370; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4371; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4372; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4373; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4374; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4375; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4376; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4377; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4378; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4379; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4380; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4381; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4382; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4383; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4384; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4385; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4386; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4387; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4388; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4389; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4390; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4391; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4392; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4393; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4394; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4395; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4396; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4397; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4398; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4399; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4400; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4401; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4402; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4403; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4404; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4405; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4406; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4407; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4408; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4409; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4410; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4411; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4412; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4413; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4414; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4415; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4416; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4417; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4418; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4419; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4420; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4421; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4422; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4423; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4424; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4425; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4426; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4427; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4428; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4429; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4430; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4431; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4432; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4433; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4434; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4435; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4436; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4437; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4438; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4439; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4440; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4441; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4442; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4443; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4444; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4445; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4446; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4447; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4448; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4449; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4450; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4451; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4452; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4453; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4454; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4455; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4456; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4457; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4458; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4459; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4460; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4461; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4462; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4463; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4464; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4465; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4466; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4467; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4468; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4469; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4470; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4471; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4472; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4473; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4474; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4475; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4476; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4477; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4478; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4479; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4480; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4481; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4482; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4483; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4484; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4485; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4486; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4487; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4488; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4489; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4490; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4491; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4492; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4493; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4494; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4495; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4496; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4497; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4498; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4499; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4500; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4501; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4502; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4503; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4504; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4505; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4506; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4507; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4508; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4509; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4510; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4511; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4512; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4513; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4514; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4515; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4516; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4517; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4518; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4519; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4520; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4521; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4522; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4523; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4524; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4525; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4526; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4527; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4528; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4529; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4530; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4531; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4532; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4533; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4534; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4535; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4536; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4537; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4538; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4539; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4540; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4541; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4542; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4543; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4544; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4545; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4546; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4547; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4548; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4549; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4550; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4551; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4552; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4553; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4554; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4555; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4556; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4557; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4558; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4559; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4560; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4561; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4562; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4563; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4564; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4565; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4566; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4567; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4568; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4569; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4570; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4571; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4572; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4573; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4574; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4575; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4576; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4577; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4578; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4579; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4580; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4581; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4582; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4583; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4584; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4585; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4586; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4587; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4588; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4589; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4590; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4591; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4592; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4593; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4594; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4595; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4596; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4597; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4598; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4599; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4600; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4601; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4602; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4603; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4604; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4605; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4606; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4607; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4608; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4609; // @[Cat.scala 30:58:@2094.4]
  wire [15:0] _T_571; // @[Cat.scala 30:58:@2094.4]
  wire [7:0] _GEN_4610; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4611; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4612; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4613; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4614; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4615; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4616; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4617; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4618; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4619; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4620; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4621; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4622; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4623; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4624; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4625; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4626; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4627; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4628; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4629; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4630; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4631; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4632; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4633; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4634; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4635; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4636; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4637; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4638; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4639; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4640; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4641; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4642; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4643; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4644; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4645; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4646; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4647; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4648; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4649; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4650; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4651; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4652; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4653; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4654; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4655; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4656; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4657; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4658; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4659; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4660; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4661; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4662; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4663; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4664; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4665; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4666; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4667; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4668; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4669; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4670; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4671; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4672; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4673; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4674; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4675; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4676; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4677; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4678; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4679; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4680; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4681; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4682; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4683; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4684; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4685; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4686; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4687; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4688; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4689; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4690; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4691; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4692; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4693; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4694; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4695; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4696; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4697; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4698; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4699; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4700; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4701; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4702; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4703; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4704; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4705; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4706; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4707; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4708; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4709; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4710; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4711; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4712; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4713; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4714; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4715; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4716; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4717; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4718; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4719; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4720; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4721; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4722; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4723; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4724; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4725; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4726; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4727; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4728; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4729; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4730; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4731; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4732; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4733; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4734; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4735; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4736; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4737; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4738; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4739; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4740; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4741; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4742; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4743; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4744; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4745; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4746; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4747; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4748; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4749; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4750; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4751; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4752; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4753; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4754; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4755; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4756; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4757; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4758; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4759; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4760; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4761; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4762; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4763; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4764; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4765; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4766; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4767; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4768; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4769; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4770; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4771; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4772; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4773; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4774; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4775; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4776; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4777; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4778; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4779; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4780; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4781; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4782; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4783; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4784; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4785; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4786; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4787; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4788; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4789; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4790; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4791; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4792; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4793; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4794; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4795; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4796; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4797; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4798; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4799; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4800; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4801; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4802; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4803; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4804; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4805; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4806; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4807; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4808; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4809; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4810; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4811; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4812; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4813; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4814; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4815; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4816; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4817; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4818; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4819; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4820; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4821; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4822; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4823; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4824; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4825; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4826; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4827; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4828; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4829; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4830; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4831; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4832; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4833; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4834; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4835; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4836; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4837; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4838; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4839; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4840; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4841; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4842; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4843; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4844; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4845; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4846; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4847; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4848; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4849; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4850; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4851; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4852; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4853; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4854; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4855; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4856; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4857; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4858; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4859; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4860; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4861; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4862; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4863; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4864; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4865; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4866; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4867; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4868; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4869; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4870; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4871; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4872; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4873; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4874; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4875; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4876; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4877; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4878; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4879; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4880; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4881; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4882; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4883; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4884; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4885; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4886; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4887; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4888; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4889; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4890; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4891; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4892; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4893; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4894; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4895; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4896; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4897; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4898; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4899; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4900; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4901; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4902; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4903; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4904; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4905; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4906; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4907; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4908; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4909; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4910; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4911; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4912; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4913; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4914; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4915; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4916; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4917; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4918; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4919; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4920; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4921; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4922; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4923; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4924; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4925; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4926; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4927; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4928; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4929; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4930; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4931; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4932; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4933; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4934; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4935; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4936; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4937; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4938; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4939; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4940; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4941; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4942; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4943; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4944; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4945; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4946; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4947; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4948; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4949; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4950; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4951; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4952; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4953; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4954; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4955; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4956; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4957; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4958; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4959; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4960; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4961; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4962; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4963; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4964; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4965; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4966; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4967; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4968; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4969; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4970; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4971; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4972; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4973; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4974; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4975; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4976; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4977; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4978; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4979; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4980; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4981; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4982; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4983; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4984; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4985; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4986; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4987; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4988; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4989; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4990; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4991; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4992; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4993; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4994; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4995; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4996; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4997; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4998; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_4999; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5000; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5001; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5002; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5003; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5004; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5005; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5006; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5007; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5008; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5009; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5010; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5011; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5012; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5013; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5014; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5015; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5016; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5017; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5018; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5019; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5020; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5021; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5022; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5023; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5024; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5025; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5026; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5027; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5028; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5029; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5030; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5031; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5032; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5033; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5034; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5035; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5036; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5037; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5038; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5039; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5040; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5041; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5042; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5043; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5044; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5045; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5046; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5047; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5048; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5049; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5050; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5051; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5052; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5053; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5054; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5055; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5056; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5057; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5058; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5059; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5060; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5061; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5062; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5063; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5064; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5065; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5066; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5067; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5068; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5069; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5070; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5071; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5072; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5073; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5074; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5075; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5076; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5077; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5078; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5079; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5080; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5081; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5082; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5083; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5084; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5085; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5086; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5087; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5088; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5089; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5090; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5091; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5092; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5093; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5094; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5095; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5096; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5097; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5098; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5099; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5100; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5101; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5102; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5103; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5104; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5105; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5106; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5107; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5108; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5109; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5110; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5111; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5112; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5113; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5114; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5115; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5116; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5117; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5118; // @[Cat.scala 30:58:@2095.4]
  wire [7:0] _GEN_5119; // @[Cat.scala 30:58:@2095.4]
  wire [15:0] _T_572; // @[Cat.scala 30:58:@2095.4]
  wire [31:0] x4; // @[Cat.scala 30:58:@2096.4]
  wire [63:0] _T_573; // @[Cat.scala 30:58:@2097.4]
  wire [63:0] _T_574; // @[Cat.scala 30:58:@2098.4]
  wire [127:0] _T_575; // @[Cat.scala 30:58:@2099.4]
  assign _T_522 = io_addr[7:0]; // @[sbox.scala 46:24:@2061.4]
  assign _T_524 = io_addr[15:8]; // @[sbox.scala 47:24:@2062.4]
  assign _T_526 = io_addr[23:16]; // @[sbox.scala 48:24:@2063.4]
  assign _T_528 = io_addr[31:24]; // @[sbox.scala 49:24:@2064.4]
  assign _GEN_20 = 8'h1 == _T_524 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_21 = 8'h2 == _T_524 ? 8'h77 : _GEN_20; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_22 = 8'h3 == _T_524 ? 8'h7b : _GEN_21; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_23 = 8'h4 == _T_524 ? 8'hf2 : _GEN_22; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_24 = 8'h5 == _T_524 ? 8'h6b : _GEN_23; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_25 = 8'h6 == _T_524 ? 8'h6f : _GEN_24; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_26 = 8'h7 == _T_524 ? 8'hc5 : _GEN_25; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_27 = 8'h8 == _T_524 ? 8'h30 : _GEN_26; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_28 = 8'h9 == _T_524 ? 8'h1 : _GEN_27; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_29 = 8'ha == _T_524 ? 8'h67 : _GEN_28; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_30 = 8'hb == _T_524 ? 8'h2b : _GEN_29; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_31 = 8'hc == _T_524 ? 8'hfe : _GEN_30; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_32 = 8'hd == _T_524 ? 8'hd7 : _GEN_31; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_33 = 8'he == _T_524 ? 8'hab : _GEN_32; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_34 = 8'hf == _T_524 ? 8'h76 : _GEN_33; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_35 = 8'h10 == _T_524 ? 8'hca : _GEN_34; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_36 = 8'h11 == _T_524 ? 8'h82 : _GEN_35; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_37 = 8'h12 == _T_524 ? 8'hc9 : _GEN_36; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_38 = 8'h13 == _T_524 ? 8'h7d : _GEN_37; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_39 = 8'h14 == _T_524 ? 8'hfa : _GEN_38; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_40 = 8'h15 == _T_524 ? 8'h59 : _GEN_39; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_41 = 8'h16 == _T_524 ? 8'h47 : _GEN_40; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_42 = 8'h17 == _T_524 ? 8'hf0 : _GEN_41; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_43 = 8'h18 == _T_524 ? 8'had : _GEN_42; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_44 = 8'h19 == _T_524 ? 8'hd4 : _GEN_43; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_45 = 8'h1a == _T_524 ? 8'ha2 : _GEN_44; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_46 = 8'h1b == _T_524 ? 8'haf : _GEN_45; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_47 = 8'h1c == _T_524 ? 8'h9c : _GEN_46; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_48 = 8'h1d == _T_524 ? 8'ha4 : _GEN_47; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_49 = 8'h1e == _T_524 ? 8'h72 : _GEN_48; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_50 = 8'h1f == _T_524 ? 8'hc0 : _GEN_49; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_51 = 8'h20 == _T_524 ? 8'hb7 : _GEN_50; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_52 = 8'h21 == _T_524 ? 8'hfd : _GEN_51; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_53 = 8'h22 == _T_524 ? 8'h93 : _GEN_52; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_54 = 8'h23 == _T_524 ? 8'h26 : _GEN_53; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_55 = 8'h24 == _T_524 ? 8'h36 : _GEN_54; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_56 = 8'h25 == _T_524 ? 8'h3f : _GEN_55; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_57 = 8'h26 == _T_524 ? 8'hf7 : _GEN_56; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_58 = 8'h27 == _T_524 ? 8'hcc : _GEN_57; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_59 = 8'h28 == _T_524 ? 8'h34 : _GEN_58; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_60 = 8'h29 == _T_524 ? 8'ha5 : _GEN_59; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_61 = 8'h2a == _T_524 ? 8'he5 : _GEN_60; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_62 = 8'h2b == _T_524 ? 8'hf1 : _GEN_61; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_63 = 8'h2c == _T_524 ? 8'h71 : _GEN_62; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_64 = 8'h2d == _T_524 ? 8'hd8 : _GEN_63; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_65 = 8'h2e == _T_524 ? 8'h31 : _GEN_64; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_66 = 8'h2f == _T_524 ? 8'h15 : _GEN_65; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_67 = 8'h30 == _T_524 ? 8'h4 : _GEN_66; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_68 = 8'h31 == _T_524 ? 8'hc7 : _GEN_67; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_69 = 8'h32 == _T_524 ? 8'h23 : _GEN_68; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_70 = 8'h33 == _T_524 ? 8'hc3 : _GEN_69; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_71 = 8'h34 == _T_524 ? 8'h18 : _GEN_70; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_72 = 8'h35 == _T_524 ? 8'h96 : _GEN_71; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_73 = 8'h36 == _T_524 ? 8'h5 : _GEN_72; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_74 = 8'h37 == _T_524 ? 8'h9a : _GEN_73; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_75 = 8'h38 == _T_524 ? 8'h7 : _GEN_74; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_76 = 8'h39 == _T_524 ? 8'h12 : _GEN_75; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_77 = 8'h3a == _T_524 ? 8'h80 : _GEN_76; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_78 = 8'h3b == _T_524 ? 8'he2 : _GEN_77; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_79 = 8'h3c == _T_524 ? 8'heb : _GEN_78; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_80 = 8'h3d == _T_524 ? 8'h27 : _GEN_79; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_81 = 8'h3e == _T_524 ? 8'hb2 : _GEN_80; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_82 = 8'h3f == _T_524 ? 8'h75 : _GEN_81; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_83 = 8'h40 == _T_524 ? 8'h9 : _GEN_82; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_84 = 8'h41 == _T_524 ? 8'h83 : _GEN_83; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_85 = 8'h42 == _T_524 ? 8'h2c : _GEN_84; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_86 = 8'h43 == _T_524 ? 8'h1a : _GEN_85; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_87 = 8'h44 == _T_524 ? 8'h1b : _GEN_86; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_88 = 8'h45 == _T_524 ? 8'h6e : _GEN_87; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_89 = 8'h46 == _T_524 ? 8'h5a : _GEN_88; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_90 = 8'h47 == _T_524 ? 8'ha0 : _GEN_89; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_91 = 8'h48 == _T_524 ? 8'h52 : _GEN_90; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_92 = 8'h49 == _T_524 ? 8'h3b : _GEN_91; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_93 = 8'h4a == _T_524 ? 8'hd6 : _GEN_92; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_94 = 8'h4b == _T_524 ? 8'hb3 : _GEN_93; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_95 = 8'h4c == _T_524 ? 8'h29 : _GEN_94; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_96 = 8'h4d == _T_524 ? 8'he3 : _GEN_95; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_97 = 8'h4e == _T_524 ? 8'h2f : _GEN_96; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_98 = 8'h4f == _T_524 ? 8'h84 : _GEN_97; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_99 = 8'h50 == _T_524 ? 8'h53 : _GEN_98; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_100 = 8'h51 == _T_524 ? 8'hd1 : _GEN_99; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_101 = 8'h52 == _T_524 ? 8'h0 : _GEN_100; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_102 = 8'h53 == _T_524 ? 8'hed : _GEN_101; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_103 = 8'h54 == _T_524 ? 8'h20 : _GEN_102; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_104 = 8'h55 == _T_524 ? 8'hfc : _GEN_103; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_105 = 8'h56 == _T_524 ? 8'hb1 : _GEN_104; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_106 = 8'h57 == _T_524 ? 8'h5b : _GEN_105; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_107 = 8'h58 == _T_524 ? 8'h6a : _GEN_106; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_108 = 8'h59 == _T_524 ? 8'hcb : _GEN_107; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_109 = 8'h5a == _T_524 ? 8'hbe : _GEN_108; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_110 = 8'h5b == _T_524 ? 8'h39 : _GEN_109; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_111 = 8'h5c == _T_524 ? 8'h4a : _GEN_110; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_112 = 8'h5d == _T_524 ? 8'h4c : _GEN_111; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_113 = 8'h5e == _T_524 ? 8'h58 : _GEN_112; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_114 = 8'h5f == _T_524 ? 8'hcf : _GEN_113; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_115 = 8'h60 == _T_524 ? 8'hd0 : _GEN_114; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_116 = 8'h61 == _T_524 ? 8'hef : _GEN_115; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_117 = 8'h62 == _T_524 ? 8'haa : _GEN_116; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_118 = 8'h63 == _T_524 ? 8'hfb : _GEN_117; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_119 = 8'h64 == _T_524 ? 8'h43 : _GEN_118; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_120 = 8'h65 == _T_524 ? 8'h4d : _GEN_119; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_121 = 8'h66 == _T_524 ? 8'h33 : _GEN_120; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_122 = 8'h67 == _T_524 ? 8'h85 : _GEN_121; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_123 = 8'h68 == _T_524 ? 8'h45 : _GEN_122; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_124 = 8'h69 == _T_524 ? 8'hf9 : _GEN_123; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_125 = 8'h6a == _T_524 ? 8'h2 : _GEN_124; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_126 = 8'h6b == _T_524 ? 8'h7f : _GEN_125; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_127 = 8'h6c == _T_524 ? 8'h50 : _GEN_126; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_128 = 8'h6d == _T_524 ? 8'h3c : _GEN_127; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_129 = 8'h6e == _T_524 ? 8'h9f : _GEN_128; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_130 = 8'h6f == _T_524 ? 8'ha8 : _GEN_129; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_131 = 8'h70 == _T_524 ? 8'h51 : _GEN_130; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_132 = 8'h71 == _T_524 ? 8'ha3 : _GEN_131; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_133 = 8'h72 == _T_524 ? 8'h40 : _GEN_132; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_134 = 8'h73 == _T_524 ? 8'h8f : _GEN_133; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_135 = 8'h74 == _T_524 ? 8'h92 : _GEN_134; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_136 = 8'h75 == _T_524 ? 8'h9d : _GEN_135; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_137 = 8'h76 == _T_524 ? 8'h38 : _GEN_136; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_138 = 8'h77 == _T_524 ? 8'hf5 : _GEN_137; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_139 = 8'h78 == _T_524 ? 8'hbc : _GEN_138; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_140 = 8'h79 == _T_524 ? 8'hb6 : _GEN_139; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_141 = 8'h7a == _T_524 ? 8'hda : _GEN_140; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_142 = 8'h7b == _T_524 ? 8'h21 : _GEN_141; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_143 = 8'h7c == _T_524 ? 8'h10 : _GEN_142; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_144 = 8'h7d == _T_524 ? 8'hff : _GEN_143; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_145 = 8'h7e == _T_524 ? 8'hf3 : _GEN_144; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_146 = 8'h7f == _T_524 ? 8'hd2 : _GEN_145; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_147 = 8'h80 == _T_524 ? 8'hcd : _GEN_146; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_148 = 8'h81 == _T_524 ? 8'hc : _GEN_147; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_149 = 8'h82 == _T_524 ? 8'h13 : _GEN_148; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_150 = 8'h83 == _T_524 ? 8'hec : _GEN_149; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_151 = 8'h84 == _T_524 ? 8'h5f : _GEN_150; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_152 = 8'h85 == _T_524 ? 8'h97 : _GEN_151; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_153 = 8'h86 == _T_524 ? 8'h44 : _GEN_152; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_154 = 8'h87 == _T_524 ? 8'h17 : _GEN_153; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_155 = 8'h88 == _T_524 ? 8'hc4 : _GEN_154; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_156 = 8'h89 == _T_524 ? 8'ha7 : _GEN_155; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_157 = 8'h8a == _T_524 ? 8'h7e : _GEN_156; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_158 = 8'h8b == _T_524 ? 8'h3d : _GEN_157; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_159 = 8'h8c == _T_524 ? 8'h64 : _GEN_158; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_160 = 8'h8d == _T_524 ? 8'h5d : _GEN_159; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_161 = 8'h8e == _T_524 ? 8'h19 : _GEN_160; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_162 = 8'h8f == _T_524 ? 8'h73 : _GEN_161; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_163 = 8'h90 == _T_524 ? 8'h60 : _GEN_162; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_164 = 8'h91 == _T_524 ? 8'h81 : _GEN_163; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_165 = 8'h92 == _T_524 ? 8'h4f : _GEN_164; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_166 = 8'h93 == _T_524 ? 8'hdc : _GEN_165; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_167 = 8'h94 == _T_524 ? 8'h22 : _GEN_166; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_168 = 8'h95 == _T_524 ? 8'h2a : _GEN_167; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_169 = 8'h96 == _T_524 ? 8'h90 : _GEN_168; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_170 = 8'h97 == _T_524 ? 8'h88 : _GEN_169; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_171 = 8'h98 == _T_524 ? 8'h46 : _GEN_170; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_172 = 8'h99 == _T_524 ? 8'hee : _GEN_171; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_173 = 8'h9a == _T_524 ? 8'hb8 : _GEN_172; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_174 = 8'h9b == _T_524 ? 8'h14 : _GEN_173; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_175 = 8'h9c == _T_524 ? 8'hde : _GEN_174; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_176 = 8'h9d == _T_524 ? 8'h5e : _GEN_175; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_177 = 8'h9e == _T_524 ? 8'hb : _GEN_176; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_178 = 8'h9f == _T_524 ? 8'hdb : _GEN_177; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_179 = 8'ha0 == _T_524 ? 8'he0 : _GEN_178; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_180 = 8'ha1 == _T_524 ? 8'h32 : _GEN_179; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_181 = 8'ha2 == _T_524 ? 8'h3a : _GEN_180; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_182 = 8'ha3 == _T_524 ? 8'ha : _GEN_181; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_183 = 8'ha4 == _T_524 ? 8'h49 : _GEN_182; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_184 = 8'ha5 == _T_524 ? 8'h6 : _GEN_183; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_185 = 8'ha6 == _T_524 ? 8'h24 : _GEN_184; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_186 = 8'ha7 == _T_524 ? 8'h5c : _GEN_185; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_187 = 8'ha8 == _T_524 ? 8'hc2 : _GEN_186; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_188 = 8'ha9 == _T_524 ? 8'hd3 : _GEN_187; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_189 = 8'haa == _T_524 ? 8'hac : _GEN_188; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_190 = 8'hab == _T_524 ? 8'h62 : _GEN_189; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_191 = 8'hac == _T_524 ? 8'h91 : _GEN_190; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_192 = 8'had == _T_524 ? 8'h95 : _GEN_191; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_193 = 8'hae == _T_524 ? 8'he4 : _GEN_192; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_194 = 8'haf == _T_524 ? 8'h79 : _GEN_193; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_195 = 8'hb0 == _T_524 ? 8'he7 : _GEN_194; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_196 = 8'hb1 == _T_524 ? 8'hc8 : _GEN_195; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_197 = 8'hb2 == _T_524 ? 8'h37 : _GEN_196; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_198 = 8'hb3 == _T_524 ? 8'h6d : _GEN_197; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_199 = 8'hb4 == _T_524 ? 8'h8d : _GEN_198; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_200 = 8'hb5 == _T_524 ? 8'hd5 : _GEN_199; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_201 = 8'hb6 == _T_524 ? 8'h4e : _GEN_200; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_202 = 8'hb7 == _T_524 ? 8'ha9 : _GEN_201; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_203 = 8'hb8 == _T_524 ? 8'h6c : _GEN_202; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_204 = 8'hb9 == _T_524 ? 8'h56 : _GEN_203; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_205 = 8'hba == _T_524 ? 8'hf4 : _GEN_204; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_206 = 8'hbb == _T_524 ? 8'hea : _GEN_205; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_207 = 8'hbc == _T_524 ? 8'h65 : _GEN_206; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_208 = 8'hbd == _T_524 ? 8'h7a : _GEN_207; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_209 = 8'hbe == _T_524 ? 8'hae : _GEN_208; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_210 = 8'hbf == _T_524 ? 8'h8 : _GEN_209; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_211 = 8'hc0 == _T_524 ? 8'hba : _GEN_210; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_212 = 8'hc1 == _T_524 ? 8'h78 : _GEN_211; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_213 = 8'hc2 == _T_524 ? 8'h25 : _GEN_212; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_214 = 8'hc3 == _T_524 ? 8'h2e : _GEN_213; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_215 = 8'hc4 == _T_524 ? 8'h1c : _GEN_214; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_216 = 8'hc5 == _T_524 ? 8'ha6 : _GEN_215; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_217 = 8'hc6 == _T_524 ? 8'hb4 : _GEN_216; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_218 = 8'hc7 == _T_524 ? 8'hc6 : _GEN_217; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_219 = 8'hc8 == _T_524 ? 8'he8 : _GEN_218; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_220 = 8'hc9 == _T_524 ? 8'hdd : _GEN_219; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_221 = 8'hca == _T_524 ? 8'h74 : _GEN_220; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_222 = 8'hcb == _T_524 ? 8'h1f : _GEN_221; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_223 = 8'hcc == _T_524 ? 8'h4b : _GEN_222; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_224 = 8'hcd == _T_524 ? 8'hbd : _GEN_223; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_225 = 8'hce == _T_524 ? 8'h8b : _GEN_224; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_226 = 8'hcf == _T_524 ? 8'h8a : _GEN_225; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_227 = 8'hd0 == _T_524 ? 8'h70 : _GEN_226; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_228 = 8'hd1 == _T_524 ? 8'h3e : _GEN_227; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_229 = 8'hd2 == _T_524 ? 8'hb5 : _GEN_228; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_230 = 8'hd3 == _T_524 ? 8'h66 : _GEN_229; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_231 = 8'hd4 == _T_524 ? 8'h48 : _GEN_230; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_232 = 8'hd5 == _T_524 ? 8'h3 : _GEN_231; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_233 = 8'hd6 == _T_524 ? 8'hf6 : _GEN_232; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_234 = 8'hd7 == _T_524 ? 8'he : _GEN_233; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_235 = 8'hd8 == _T_524 ? 8'h61 : _GEN_234; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_236 = 8'hd9 == _T_524 ? 8'h35 : _GEN_235; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_237 = 8'hda == _T_524 ? 8'h57 : _GEN_236; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_238 = 8'hdb == _T_524 ? 8'hb9 : _GEN_237; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_239 = 8'hdc == _T_524 ? 8'h86 : _GEN_238; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_240 = 8'hdd == _T_524 ? 8'hc1 : _GEN_239; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_241 = 8'hde == _T_524 ? 8'h1d : _GEN_240; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_242 = 8'hdf == _T_524 ? 8'h9e : _GEN_241; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_243 = 8'he0 == _T_524 ? 8'he1 : _GEN_242; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_244 = 8'he1 == _T_524 ? 8'hf8 : _GEN_243; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_245 = 8'he2 == _T_524 ? 8'h98 : _GEN_244; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_246 = 8'he3 == _T_524 ? 8'h11 : _GEN_245; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_247 = 8'he4 == _T_524 ? 8'h69 : _GEN_246; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_248 = 8'he5 == _T_524 ? 8'hd9 : _GEN_247; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_249 = 8'he6 == _T_524 ? 8'h8e : _GEN_248; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_250 = 8'he7 == _T_524 ? 8'h94 : _GEN_249; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_251 = 8'he8 == _T_524 ? 8'h9b : _GEN_250; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_252 = 8'he9 == _T_524 ? 8'h1e : _GEN_251; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_253 = 8'hea == _T_524 ? 8'h87 : _GEN_252; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_254 = 8'heb == _T_524 ? 8'he9 : _GEN_253; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_255 = 8'hec == _T_524 ? 8'hce : _GEN_254; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_256 = 8'hed == _T_524 ? 8'h55 : _GEN_255; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_257 = 8'hee == _T_524 ? 8'h28 : _GEN_256; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_258 = 8'hef == _T_524 ? 8'hdf : _GEN_257; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_259 = 8'hf0 == _T_524 ? 8'h8c : _GEN_258; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_260 = 8'hf1 == _T_524 ? 8'ha1 : _GEN_259; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_261 = 8'hf2 == _T_524 ? 8'h89 : _GEN_260; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_262 = 8'hf3 == _T_524 ? 8'hd : _GEN_261; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_263 = 8'hf4 == _T_524 ? 8'hbf : _GEN_262; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_264 = 8'hf5 == _T_524 ? 8'he6 : _GEN_263; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_265 = 8'hf6 == _T_524 ? 8'h42 : _GEN_264; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_266 = 8'hf7 == _T_524 ? 8'h68 : _GEN_265; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_267 = 8'hf8 == _T_524 ? 8'h41 : _GEN_266; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_268 = 8'hf9 == _T_524 ? 8'h99 : _GEN_267; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_269 = 8'hfa == _T_524 ? 8'h2d : _GEN_268; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_270 = 8'hfb == _T_524 ? 8'hf : _GEN_269; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_271 = 8'hfc == _T_524 ? 8'hb0 : _GEN_270; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_272 = 8'hfd == _T_524 ? 8'h54 : _GEN_271; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_273 = 8'hfe == _T_524 ? 8'hbb : _GEN_272; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_274 = 8'hff == _T_524 ? 8'h16 : _GEN_273; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_275 = 8'h1 == _T_522 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_276 = 8'h2 == _T_522 ? 8'h77 : _GEN_275; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_277 = 8'h3 == _T_522 ? 8'h7b : _GEN_276; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_278 = 8'h4 == _T_522 ? 8'hf2 : _GEN_277; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_279 = 8'h5 == _T_522 ? 8'h6b : _GEN_278; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_280 = 8'h6 == _T_522 ? 8'h6f : _GEN_279; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_281 = 8'h7 == _T_522 ? 8'hc5 : _GEN_280; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_282 = 8'h8 == _T_522 ? 8'h30 : _GEN_281; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_283 = 8'h9 == _T_522 ? 8'h1 : _GEN_282; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_284 = 8'ha == _T_522 ? 8'h67 : _GEN_283; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_285 = 8'hb == _T_522 ? 8'h2b : _GEN_284; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_286 = 8'hc == _T_522 ? 8'hfe : _GEN_285; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_287 = 8'hd == _T_522 ? 8'hd7 : _GEN_286; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_288 = 8'he == _T_522 ? 8'hab : _GEN_287; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_289 = 8'hf == _T_522 ? 8'h76 : _GEN_288; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_290 = 8'h10 == _T_522 ? 8'hca : _GEN_289; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_291 = 8'h11 == _T_522 ? 8'h82 : _GEN_290; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_292 = 8'h12 == _T_522 ? 8'hc9 : _GEN_291; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_293 = 8'h13 == _T_522 ? 8'h7d : _GEN_292; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_294 = 8'h14 == _T_522 ? 8'hfa : _GEN_293; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_295 = 8'h15 == _T_522 ? 8'h59 : _GEN_294; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_296 = 8'h16 == _T_522 ? 8'h47 : _GEN_295; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_297 = 8'h17 == _T_522 ? 8'hf0 : _GEN_296; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_298 = 8'h18 == _T_522 ? 8'had : _GEN_297; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_299 = 8'h19 == _T_522 ? 8'hd4 : _GEN_298; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_300 = 8'h1a == _T_522 ? 8'ha2 : _GEN_299; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_301 = 8'h1b == _T_522 ? 8'haf : _GEN_300; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_302 = 8'h1c == _T_522 ? 8'h9c : _GEN_301; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_303 = 8'h1d == _T_522 ? 8'ha4 : _GEN_302; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_304 = 8'h1e == _T_522 ? 8'h72 : _GEN_303; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_305 = 8'h1f == _T_522 ? 8'hc0 : _GEN_304; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_306 = 8'h20 == _T_522 ? 8'hb7 : _GEN_305; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_307 = 8'h21 == _T_522 ? 8'hfd : _GEN_306; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_308 = 8'h22 == _T_522 ? 8'h93 : _GEN_307; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_309 = 8'h23 == _T_522 ? 8'h26 : _GEN_308; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_310 = 8'h24 == _T_522 ? 8'h36 : _GEN_309; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_311 = 8'h25 == _T_522 ? 8'h3f : _GEN_310; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_312 = 8'h26 == _T_522 ? 8'hf7 : _GEN_311; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_313 = 8'h27 == _T_522 ? 8'hcc : _GEN_312; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_314 = 8'h28 == _T_522 ? 8'h34 : _GEN_313; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_315 = 8'h29 == _T_522 ? 8'ha5 : _GEN_314; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_316 = 8'h2a == _T_522 ? 8'he5 : _GEN_315; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_317 = 8'h2b == _T_522 ? 8'hf1 : _GEN_316; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_318 = 8'h2c == _T_522 ? 8'h71 : _GEN_317; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_319 = 8'h2d == _T_522 ? 8'hd8 : _GEN_318; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_320 = 8'h2e == _T_522 ? 8'h31 : _GEN_319; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_321 = 8'h2f == _T_522 ? 8'h15 : _GEN_320; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_322 = 8'h30 == _T_522 ? 8'h4 : _GEN_321; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_323 = 8'h31 == _T_522 ? 8'hc7 : _GEN_322; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_324 = 8'h32 == _T_522 ? 8'h23 : _GEN_323; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_325 = 8'h33 == _T_522 ? 8'hc3 : _GEN_324; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_326 = 8'h34 == _T_522 ? 8'h18 : _GEN_325; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_327 = 8'h35 == _T_522 ? 8'h96 : _GEN_326; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_328 = 8'h36 == _T_522 ? 8'h5 : _GEN_327; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_329 = 8'h37 == _T_522 ? 8'h9a : _GEN_328; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_330 = 8'h38 == _T_522 ? 8'h7 : _GEN_329; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_331 = 8'h39 == _T_522 ? 8'h12 : _GEN_330; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_332 = 8'h3a == _T_522 ? 8'h80 : _GEN_331; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_333 = 8'h3b == _T_522 ? 8'he2 : _GEN_332; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_334 = 8'h3c == _T_522 ? 8'heb : _GEN_333; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_335 = 8'h3d == _T_522 ? 8'h27 : _GEN_334; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_336 = 8'h3e == _T_522 ? 8'hb2 : _GEN_335; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_337 = 8'h3f == _T_522 ? 8'h75 : _GEN_336; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_338 = 8'h40 == _T_522 ? 8'h9 : _GEN_337; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_339 = 8'h41 == _T_522 ? 8'h83 : _GEN_338; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_340 = 8'h42 == _T_522 ? 8'h2c : _GEN_339; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_341 = 8'h43 == _T_522 ? 8'h1a : _GEN_340; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_342 = 8'h44 == _T_522 ? 8'h1b : _GEN_341; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_343 = 8'h45 == _T_522 ? 8'h6e : _GEN_342; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_344 = 8'h46 == _T_522 ? 8'h5a : _GEN_343; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_345 = 8'h47 == _T_522 ? 8'ha0 : _GEN_344; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_346 = 8'h48 == _T_522 ? 8'h52 : _GEN_345; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_347 = 8'h49 == _T_522 ? 8'h3b : _GEN_346; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_348 = 8'h4a == _T_522 ? 8'hd6 : _GEN_347; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_349 = 8'h4b == _T_522 ? 8'hb3 : _GEN_348; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_350 = 8'h4c == _T_522 ? 8'h29 : _GEN_349; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_351 = 8'h4d == _T_522 ? 8'he3 : _GEN_350; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_352 = 8'h4e == _T_522 ? 8'h2f : _GEN_351; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_353 = 8'h4f == _T_522 ? 8'h84 : _GEN_352; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_354 = 8'h50 == _T_522 ? 8'h53 : _GEN_353; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_355 = 8'h51 == _T_522 ? 8'hd1 : _GEN_354; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_356 = 8'h52 == _T_522 ? 8'h0 : _GEN_355; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_357 = 8'h53 == _T_522 ? 8'hed : _GEN_356; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_358 = 8'h54 == _T_522 ? 8'h20 : _GEN_357; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_359 = 8'h55 == _T_522 ? 8'hfc : _GEN_358; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_360 = 8'h56 == _T_522 ? 8'hb1 : _GEN_359; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_361 = 8'h57 == _T_522 ? 8'h5b : _GEN_360; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_362 = 8'h58 == _T_522 ? 8'h6a : _GEN_361; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_363 = 8'h59 == _T_522 ? 8'hcb : _GEN_362; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_364 = 8'h5a == _T_522 ? 8'hbe : _GEN_363; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_365 = 8'h5b == _T_522 ? 8'h39 : _GEN_364; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_366 = 8'h5c == _T_522 ? 8'h4a : _GEN_365; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_367 = 8'h5d == _T_522 ? 8'h4c : _GEN_366; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_368 = 8'h5e == _T_522 ? 8'h58 : _GEN_367; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_369 = 8'h5f == _T_522 ? 8'hcf : _GEN_368; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_370 = 8'h60 == _T_522 ? 8'hd0 : _GEN_369; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_371 = 8'h61 == _T_522 ? 8'hef : _GEN_370; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_372 = 8'h62 == _T_522 ? 8'haa : _GEN_371; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_373 = 8'h63 == _T_522 ? 8'hfb : _GEN_372; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_374 = 8'h64 == _T_522 ? 8'h43 : _GEN_373; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_375 = 8'h65 == _T_522 ? 8'h4d : _GEN_374; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_376 = 8'h66 == _T_522 ? 8'h33 : _GEN_375; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_377 = 8'h67 == _T_522 ? 8'h85 : _GEN_376; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_378 = 8'h68 == _T_522 ? 8'h45 : _GEN_377; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_379 = 8'h69 == _T_522 ? 8'hf9 : _GEN_378; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_380 = 8'h6a == _T_522 ? 8'h2 : _GEN_379; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_381 = 8'h6b == _T_522 ? 8'h7f : _GEN_380; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_382 = 8'h6c == _T_522 ? 8'h50 : _GEN_381; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_383 = 8'h6d == _T_522 ? 8'h3c : _GEN_382; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_384 = 8'h6e == _T_522 ? 8'h9f : _GEN_383; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_385 = 8'h6f == _T_522 ? 8'ha8 : _GEN_384; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_386 = 8'h70 == _T_522 ? 8'h51 : _GEN_385; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_387 = 8'h71 == _T_522 ? 8'ha3 : _GEN_386; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_388 = 8'h72 == _T_522 ? 8'h40 : _GEN_387; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_389 = 8'h73 == _T_522 ? 8'h8f : _GEN_388; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_390 = 8'h74 == _T_522 ? 8'h92 : _GEN_389; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_391 = 8'h75 == _T_522 ? 8'h9d : _GEN_390; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_392 = 8'h76 == _T_522 ? 8'h38 : _GEN_391; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_393 = 8'h77 == _T_522 ? 8'hf5 : _GEN_392; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_394 = 8'h78 == _T_522 ? 8'hbc : _GEN_393; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_395 = 8'h79 == _T_522 ? 8'hb6 : _GEN_394; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_396 = 8'h7a == _T_522 ? 8'hda : _GEN_395; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_397 = 8'h7b == _T_522 ? 8'h21 : _GEN_396; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_398 = 8'h7c == _T_522 ? 8'h10 : _GEN_397; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_399 = 8'h7d == _T_522 ? 8'hff : _GEN_398; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_400 = 8'h7e == _T_522 ? 8'hf3 : _GEN_399; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_401 = 8'h7f == _T_522 ? 8'hd2 : _GEN_400; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_402 = 8'h80 == _T_522 ? 8'hcd : _GEN_401; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_403 = 8'h81 == _T_522 ? 8'hc : _GEN_402; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_404 = 8'h82 == _T_522 ? 8'h13 : _GEN_403; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_405 = 8'h83 == _T_522 ? 8'hec : _GEN_404; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_406 = 8'h84 == _T_522 ? 8'h5f : _GEN_405; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_407 = 8'h85 == _T_522 ? 8'h97 : _GEN_406; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_408 = 8'h86 == _T_522 ? 8'h44 : _GEN_407; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_409 = 8'h87 == _T_522 ? 8'h17 : _GEN_408; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_410 = 8'h88 == _T_522 ? 8'hc4 : _GEN_409; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_411 = 8'h89 == _T_522 ? 8'ha7 : _GEN_410; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_412 = 8'h8a == _T_522 ? 8'h7e : _GEN_411; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_413 = 8'h8b == _T_522 ? 8'h3d : _GEN_412; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_414 = 8'h8c == _T_522 ? 8'h64 : _GEN_413; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_415 = 8'h8d == _T_522 ? 8'h5d : _GEN_414; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_416 = 8'h8e == _T_522 ? 8'h19 : _GEN_415; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_417 = 8'h8f == _T_522 ? 8'h73 : _GEN_416; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_418 = 8'h90 == _T_522 ? 8'h60 : _GEN_417; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_419 = 8'h91 == _T_522 ? 8'h81 : _GEN_418; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_420 = 8'h92 == _T_522 ? 8'h4f : _GEN_419; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_421 = 8'h93 == _T_522 ? 8'hdc : _GEN_420; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_422 = 8'h94 == _T_522 ? 8'h22 : _GEN_421; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_423 = 8'h95 == _T_522 ? 8'h2a : _GEN_422; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_424 = 8'h96 == _T_522 ? 8'h90 : _GEN_423; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_425 = 8'h97 == _T_522 ? 8'h88 : _GEN_424; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_426 = 8'h98 == _T_522 ? 8'h46 : _GEN_425; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_427 = 8'h99 == _T_522 ? 8'hee : _GEN_426; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_428 = 8'h9a == _T_522 ? 8'hb8 : _GEN_427; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_429 = 8'h9b == _T_522 ? 8'h14 : _GEN_428; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_430 = 8'h9c == _T_522 ? 8'hde : _GEN_429; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_431 = 8'h9d == _T_522 ? 8'h5e : _GEN_430; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_432 = 8'h9e == _T_522 ? 8'hb : _GEN_431; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_433 = 8'h9f == _T_522 ? 8'hdb : _GEN_432; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_434 = 8'ha0 == _T_522 ? 8'he0 : _GEN_433; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_435 = 8'ha1 == _T_522 ? 8'h32 : _GEN_434; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_436 = 8'ha2 == _T_522 ? 8'h3a : _GEN_435; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_437 = 8'ha3 == _T_522 ? 8'ha : _GEN_436; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_438 = 8'ha4 == _T_522 ? 8'h49 : _GEN_437; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_439 = 8'ha5 == _T_522 ? 8'h6 : _GEN_438; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_440 = 8'ha6 == _T_522 ? 8'h24 : _GEN_439; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_441 = 8'ha7 == _T_522 ? 8'h5c : _GEN_440; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_442 = 8'ha8 == _T_522 ? 8'hc2 : _GEN_441; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_443 = 8'ha9 == _T_522 ? 8'hd3 : _GEN_442; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_444 = 8'haa == _T_522 ? 8'hac : _GEN_443; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_445 = 8'hab == _T_522 ? 8'h62 : _GEN_444; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_446 = 8'hac == _T_522 ? 8'h91 : _GEN_445; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_447 = 8'had == _T_522 ? 8'h95 : _GEN_446; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_448 = 8'hae == _T_522 ? 8'he4 : _GEN_447; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_449 = 8'haf == _T_522 ? 8'h79 : _GEN_448; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_450 = 8'hb0 == _T_522 ? 8'he7 : _GEN_449; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_451 = 8'hb1 == _T_522 ? 8'hc8 : _GEN_450; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_452 = 8'hb2 == _T_522 ? 8'h37 : _GEN_451; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_453 = 8'hb3 == _T_522 ? 8'h6d : _GEN_452; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_454 = 8'hb4 == _T_522 ? 8'h8d : _GEN_453; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_455 = 8'hb5 == _T_522 ? 8'hd5 : _GEN_454; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_456 = 8'hb6 == _T_522 ? 8'h4e : _GEN_455; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_457 = 8'hb7 == _T_522 ? 8'ha9 : _GEN_456; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_458 = 8'hb8 == _T_522 ? 8'h6c : _GEN_457; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_459 = 8'hb9 == _T_522 ? 8'h56 : _GEN_458; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_460 = 8'hba == _T_522 ? 8'hf4 : _GEN_459; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_461 = 8'hbb == _T_522 ? 8'hea : _GEN_460; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_462 = 8'hbc == _T_522 ? 8'h65 : _GEN_461; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_463 = 8'hbd == _T_522 ? 8'h7a : _GEN_462; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_464 = 8'hbe == _T_522 ? 8'hae : _GEN_463; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_465 = 8'hbf == _T_522 ? 8'h8 : _GEN_464; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_466 = 8'hc0 == _T_522 ? 8'hba : _GEN_465; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_467 = 8'hc1 == _T_522 ? 8'h78 : _GEN_466; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_468 = 8'hc2 == _T_522 ? 8'h25 : _GEN_467; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_469 = 8'hc3 == _T_522 ? 8'h2e : _GEN_468; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_470 = 8'hc4 == _T_522 ? 8'h1c : _GEN_469; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_471 = 8'hc5 == _T_522 ? 8'ha6 : _GEN_470; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_472 = 8'hc6 == _T_522 ? 8'hb4 : _GEN_471; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_473 = 8'hc7 == _T_522 ? 8'hc6 : _GEN_472; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_474 = 8'hc8 == _T_522 ? 8'he8 : _GEN_473; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_475 = 8'hc9 == _T_522 ? 8'hdd : _GEN_474; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_476 = 8'hca == _T_522 ? 8'h74 : _GEN_475; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_477 = 8'hcb == _T_522 ? 8'h1f : _GEN_476; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_478 = 8'hcc == _T_522 ? 8'h4b : _GEN_477; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_479 = 8'hcd == _T_522 ? 8'hbd : _GEN_478; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_480 = 8'hce == _T_522 ? 8'h8b : _GEN_479; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_481 = 8'hcf == _T_522 ? 8'h8a : _GEN_480; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_482 = 8'hd0 == _T_522 ? 8'h70 : _GEN_481; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_483 = 8'hd1 == _T_522 ? 8'h3e : _GEN_482; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_484 = 8'hd2 == _T_522 ? 8'hb5 : _GEN_483; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_485 = 8'hd3 == _T_522 ? 8'h66 : _GEN_484; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_486 = 8'hd4 == _T_522 ? 8'h48 : _GEN_485; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_487 = 8'hd5 == _T_522 ? 8'h3 : _GEN_486; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_488 = 8'hd6 == _T_522 ? 8'hf6 : _GEN_487; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_489 = 8'hd7 == _T_522 ? 8'he : _GEN_488; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_490 = 8'hd8 == _T_522 ? 8'h61 : _GEN_489; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_491 = 8'hd9 == _T_522 ? 8'h35 : _GEN_490; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_492 = 8'hda == _T_522 ? 8'h57 : _GEN_491; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_493 = 8'hdb == _T_522 ? 8'hb9 : _GEN_492; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_494 = 8'hdc == _T_522 ? 8'h86 : _GEN_493; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_495 = 8'hdd == _T_522 ? 8'hc1 : _GEN_494; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_496 = 8'hde == _T_522 ? 8'h1d : _GEN_495; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_497 = 8'hdf == _T_522 ? 8'h9e : _GEN_496; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_498 = 8'he0 == _T_522 ? 8'he1 : _GEN_497; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_499 = 8'he1 == _T_522 ? 8'hf8 : _GEN_498; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_500 = 8'he2 == _T_522 ? 8'h98 : _GEN_499; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_501 = 8'he3 == _T_522 ? 8'h11 : _GEN_500; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_502 = 8'he4 == _T_522 ? 8'h69 : _GEN_501; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_503 = 8'he5 == _T_522 ? 8'hd9 : _GEN_502; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_504 = 8'he6 == _T_522 ? 8'h8e : _GEN_503; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_505 = 8'he7 == _T_522 ? 8'h94 : _GEN_504; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_506 = 8'he8 == _T_522 ? 8'h9b : _GEN_505; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_507 = 8'he9 == _T_522 ? 8'h1e : _GEN_506; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_508 = 8'hea == _T_522 ? 8'h87 : _GEN_507; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_509 = 8'heb == _T_522 ? 8'he9 : _GEN_508; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_510 = 8'hec == _T_522 ? 8'hce : _GEN_509; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_511 = 8'hed == _T_522 ? 8'h55 : _GEN_510; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_512 = 8'hee == _T_522 ? 8'h28 : _GEN_511; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_513 = 8'hef == _T_522 ? 8'hdf : _GEN_512; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_514 = 8'hf0 == _T_522 ? 8'h8c : _GEN_513; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_515 = 8'hf1 == _T_522 ? 8'ha1 : _GEN_514; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_516 = 8'hf2 == _T_522 ? 8'h89 : _GEN_515; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_517 = 8'hf3 == _T_522 ? 8'hd : _GEN_516; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_518 = 8'hf4 == _T_522 ? 8'hbf : _GEN_517; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_519 = 8'hf5 == _T_522 ? 8'he6 : _GEN_518; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_520 = 8'hf6 == _T_522 ? 8'h42 : _GEN_519; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_521 = 8'hf7 == _T_522 ? 8'h68 : _GEN_520; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_522 = 8'hf8 == _T_522 ? 8'h41 : _GEN_521; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_523 = 8'hf9 == _T_522 ? 8'h99 : _GEN_522; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_524 = 8'hfa == _T_522 ? 8'h2d : _GEN_523; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_525 = 8'hfb == _T_522 ? 8'hf : _GEN_524; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_526 = 8'hfc == _T_522 ? 8'hb0 : _GEN_525; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_527 = 8'hfd == _T_522 ? 8'h54 : _GEN_526; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_528 = 8'hfe == _T_522 ? 8'hbb : _GEN_527; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_529 = 8'hff == _T_522 ? 8'h16 : _GEN_528; // @[Cat.scala 30:58:@2065.4]
  assign _T_530 = {_GEN_274,_GEN_529}; // @[Cat.scala 30:58:@2065.4]
  assign _GEN_530 = 8'h1 == _T_528 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_531 = 8'h2 == _T_528 ? 8'h77 : _GEN_530; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_532 = 8'h3 == _T_528 ? 8'h7b : _GEN_531; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_533 = 8'h4 == _T_528 ? 8'hf2 : _GEN_532; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_534 = 8'h5 == _T_528 ? 8'h6b : _GEN_533; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_535 = 8'h6 == _T_528 ? 8'h6f : _GEN_534; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_536 = 8'h7 == _T_528 ? 8'hc5 : _GEN_535; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_537 = 8'h8 == _T_528 ? 8'h30 : _GEN_536; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_538 = 8'h9 == _T_528 ? 8'h1 : _GEN_537; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_539 = 8'ha == _T_528 ? 8'h67 : _GEN_538; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_540 = 8'hb == _T_528 ? 8'h2b : _GEN_539; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_541 = 8'hc == _T_528 ? 8'hfe : _GEN_540; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_542 = 8'hd == _T_528 ? 8'hd7 : _GEN_541; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_543 = 8'he == _T_528 ? 8'hab : _GEN_542; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_544 = 8'hf == _T_528 ? 8'h76 : _GEN_543; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_545 = 8'h10 == _T_528 ? 8'hca : _GEN_544; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_546 = 8'h11 == _T_528 ? 8'h82 : _GEN_545; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_547 = 8'h12 == _T_528 ? 8'hc9 : _GEN_546; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_548 = 8'h13 == _T_528 ? 8'h7d : _GEN_547; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_549 = 8'h14 == _T_528 ? 8'hfa : _GEN_548; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_550 = 8'h15 == _T_528 ? 8'h59 : _GEN_549; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_551 = 8'h16 == _T_528 ? 8'h47 : _GEN_550; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_552 = 8'h17 == _T_528 ? 8'hf0 : _GEN_551; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_553 = 8'h18 == _T_528 ? 8'had : _GEN_552; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_554 = 8'h19 == _T_528 ? 8'hd4 : _GEN_553; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_555 = 8'h1a == _T_528 ? 8'ha2 : _GEN_554; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_556 = 8'h1b == _T_528 ? 8'haf : _GEN_555; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_557 = 8'h1c == _T_528 ? 8'h9c : _GEN_556; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_558 = 8'h1d == _T_528 ? 8'ha4 : _GEN_557; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_559 = 8'h1e == _T_528 ? 8'h72 : _GEN_558; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_560 = 8'h1f == _T_528 ? 8'hc0 : _GEN_559; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_561 = 8'h20 == _T_528 ? 8'hb7 : _GEN_560; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_562 = 8'h21 == _T_528 ? 8'hfd : _GEN_561; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_563 = 8'h22 == _T_528 ? 8'h93 : _GEN_562; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_564 = 8'h23 == _T_528 ? 8'h26 : _GEN_563; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_565 = 8'h24 == _T_528 ? 8'h36 : _GEN_564; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_566 = 8'h25 == _T_528 ? 8'h3f : _GEN_565; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_567 = 8'h26 == _T_528 ? 8'hf7 : _GEN_566; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_568 = 8'h27 == _T_528 ? 8'hcc : _GEN_567; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_569 = 8'h28 == _T_528 ? 8'h34 : _GEN_568; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_570 = 8'h29 == _T_528 ? 8'ha5 : _GEN_569; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_571 = 8'h2a == _T_528 ? 8'he5 : _GEN_570; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_572 = 8'h2b == _T_528 ? 8'hf1 : _GEN_571; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_573 = 8'h2c == _T_528 ? 8'h71 : _GEN_572; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_574 = 8'h2d == _T_528 ? 8'hd8 : _GEN_573; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_575 = 8'h2e == _T_528 ? 8'h31 : _GEN_574; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_576 = 8'h2f == _T_528 ? 8'h15 : _GEN_575; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_577 = 8'h30 == _T_528 ? 8'h4 : _GEN_576; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_578 = 8'h31 == _T_528 ? 8'hc7 : _GEN_577; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_579 = 8'h32 == _T_528 ? 8'h23 : _GEN_578; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_580 = 8'h33 == _T_528 ? 8'hc3 : _GEN_579; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_581 = 8'h34 == _T_528 ? 8'h18 : _GEN_580; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_582 = 8'h35 == _T_528 ? 8'h96 : _GEN_581; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_583 = 8'h36 == _T_528 ? 8'h5 : _GEN_582; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_584 = 8'h37 == _T_528 ? 8'h9a : _GEN_583; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_585 = 8'h38 == _T_528 ? 8'h7 : _GEN_584; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_586 = 8'h39 == _T_528 ? 8'h12 : _GEN_585; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_587 = 8'h3a == _T_528 ? 8'h80 : _GEN_586; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_588 = 8'h3b == _T_528 ? 8'he2 : _GEN_587; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_589 = 8'h3c == _T_528 ? 8'heb : _GEN_588; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_590 = 8'h3d == _T_528 ? 8'h27 : _GEN_589; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_591 = 8'h3e == _T_528 ? 8'hb2 : _GEN_590; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_592 = 8'h3f == _T_528 ? 8'h75 : _GEN_591; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_593 = 8'h40 == _T_528 ? 8'h9 : _GEN_592; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_594 = 8'h41 == _T_528 ? 8'h83 : _GEN_593; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_595 = 8'h42 == _T_528 ? 8'h2c : _GEN_594; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_596 = 8'h43 == _T_528 ? 8'h1a : _GEN_595; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_597 = 8'h44 == _T_528 ? 8'h1b : _GEN_596; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_598 = 8'h45 == _T_528 ? 8'h6e : _GEN_597; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_599 = 8'h46 == _T_528 ? 8'h5a : _GEN_598; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_600 = 8'h47 == _T_528 ? 8'ha0 : _GEN_599; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_601 = 8'h48 == _T_528 ? 8'h52 : _GEN_600; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_602 = 8'h49 == _T_528 ? 8'h3b : _GEN_601; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_603 = 8'h4a == _T_528 ? 8'hd6 : _GEN_602; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_604 = 8'h4b == _T_528 ? 8'hb3 : _GEN_603; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_605 = 8'h4c == _T_528 ? 8'h29 : _GEN_604; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_606 = 8'h4d == _T_528 ? 8'he3 : _GEN_605; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_607 = 8'h4e == _T_528 ? 8'h2f : _GEN_606; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_608 = 8'h4f == _T_528 ? 8'h84 : _GEN_607; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_609 = 8'h50 == _T_528 ? 8'h53 : _GEN_608; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_610 = 8'h51 == _T_528 ? 8'hd1 : _GEN_609; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_611 = 8'h52 == _T_528 ? 8'h0 : _GEN_610; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_612 = 8'h53 == _T_528 ? 8'hed : _GEN_611; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_613 = 8'h54 == _T_528 ? 8'h20 : _GEN_612; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_614 = 8'h55 == _T_528 ? 8'hfc : _GEN_613; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_615 = 8'h56 == _T_528 ? 8'hb1 : _GEN_614; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_616 = 8'h57 == _T_528 ? 8'h5b : _GEN_615; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_617 = 8'h58 == _T_528 ? 8'h6a : _GEN_616; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_618 = 8'h59 == _T_528 ? 8'hcb : _GEN_617; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_619 = 8'h5a == _T_528 ? 8'hbe : _GEN_618; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_620 = 8'h5b == _T_528 ? 8'h39 : _GEN_619; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_621 = 8'h5c == _T_528 ? 8'h4a : _GEN_620; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_622 = 8'h5d == _T_528 ? 8'h4c : _GEN_621; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_623 = 8'h5e == _T_528 ? 8'h58 : _GEN_622; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_624 = 8'h5f == _T_528 ? 8'hcf : _GEN_623; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_625 = 8'h60 == _T_528 ? 8'hd0 : _GEN_624; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_626 = 8'h61 == _T_528 ? 8'hef : _GEN_625; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_627 = 8'h62 == _T_528 ? 8'haa : _GEN_626; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_628 = 8'h63 == _T_528 ? 8'hfb : _GEN_627; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_629 = 8'h64 == _T_528 ? 8'h43 : _GEN_628; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_630 = 8'h65 == _T_528 ? 8'h4d : _GEN_629; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_631 = 8'h66 == _T_528 ? 8'h33 : _GEN_630; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_632 = 8'h67 == _T_528 ? 8'h85 : _GEN_631; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_633 = 8'h68 == _T_528 ? 8'h45 : _GEN_632; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_634 = 8'h69 == _T_528 ? 8'hf9 : _GEN_633; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_635 = 8'h6a == _T_528 ? 8'h2 : _GEN_634; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_636 = 8'h6b == _T_528 ? 8'h7f : _GEN_635; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_637 = 8'h6c == _T_528 ? 8'h50 : _GEN_636; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_638 = 8'h6d == _T_528 ? 8'h3c : _GEN_637; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_639 = 8'h6e == _T_528 ? 8'h9f : _GEN_638; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_640 = 8'h6f == _T_528 ? 8'ha8 : _GEN_639; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_641 = 8'h70 == _T_528 ? 8'h51 : _GEN_640; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_642 = 8'h71 == _T_528 ? 8'ha3 : _GEN_641; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_643 = 8'h72 == _T_528 ? 8'h40 : _GEN_642; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_644 = 8'h73 == _T_528 ? 8'h8f : _GEN_643; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_645 = 8'h74 == _T_528 ? 8'h92 : _GEN_644; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_646 = 8'h75 == _T_528 ? 8'h9d : _GEN_645; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_647 = 8'h76 == _T_528 ? 8'h38 : _GEN_646; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_648 = 8'h77 == _T_528 ? 8'hf5 : _GEN_647; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_649 = 8'h78 == _T_528 ? 8'hbc : _GEN_648; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_650 = 8'h79 == _T_528 ? 8'hb6 : _GEN_649; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_651 = 8'h7a == _T_528 ? 8'hda : _GEN_650; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_652 = 8'h7b == _T_528 ? 8'h21 : _GEN_651; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_653 = 8'h7c == _T_528 ? 8'h10 : _GEN_652; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_654 = 8'h7d == _T_528 ? 8'hff : _GEN_653; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_655 = 8'h7e == _T_528 ? 8'hf3 : _GEN_654; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_656 = 8'h7f == _T_528 ? 8'hd2 : _GEN_655; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_657 = 8'h80 == _T_528 ? 8'hcd : _GEN_656; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_658 = 8'h81 == _T_528 ? 8'hc : _GEN_657; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_659 = 8'h82 == _T_528 ? 8'h13 : _GEN_658; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_660 = 8'h83 == _T_528 ? 8'hec : _GEN_659; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_661 = 8'h84 == _T_528 ? 8'h5f : _GEN_660; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_662 = 8'h85 == _T_528 ? 8'h97 : _GEN_661; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_663 = 8'h86 == _T_528 ? 8'h44 : _GEN_662; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_664 = 8'h87 == _T_528 ? 8'h17 : _GEN_663; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_665 = 8'h88 == _T_528 ? 8'hc4 : _GEN_664; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_666 = 8'h89 == _T_528 ? 8'ha7 : _GEN_665; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_667 = 8'h8a == _T_528 ? 8'h7e : _GEN_666; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_668 = 8'h8b == _T_528 ? 8'h3d : _GEN_667; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_669 = 8'h8c == _T_528 ? 8'h64 : _GEN_668; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_670 = 8'h8d == _T_528 ? 8'h5d : _GEN_669; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_671 = 8'h8e == _T_528 ? 8'h19 : _GEN_670; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_672 = 8'h8f == _T_528 ? 8'h73 : _GEN_671; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_673 = 8'h90 == _T_528 ? 8'h60 : _GEN_672; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_674 = 8'h91 == _T_528 ? 8'h81 : _GEN_673; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_675 = 8'h92 == _T_528 ? 8'h4f : _GEN_674; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_676 = 8'h93 == _T_528 ? 8'hdc : _GEN_675; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_677 = 8'h94 == _T_528 ? 8'h22 : _GEN_676; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_678 = 8'h95 == _T_528 ? 8'h2a : _GEN_677; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_679 = 8'h96 == _T_528 ? 8'h90 : _GEN_678; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_680 = 8'h97 == _T_528 ? 8'h88 : _GEN_679; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_681 = 8'h98 == _T_528 ? 8'h46 : _GEN_680; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_682 = 8'h99 == _T_528 ? 8'hee : _GEN_681; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_683 = 8'h9a == _T_528 ? 8'hb8 : _GEN_682; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_684 = 8'h9b == _T_528 ? 8'h14 : _GEN_683; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_685 = 8'h9c == _T_528 ? 8'hde : _GEN_684; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_686 = 8'h9d == _T_528 ? 8'h5e : _GEN_685; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_687 = 8'h9e == _T_528 ? 8'hb : _GEN_686; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_688 = 8'h9f == _T_528 ? 8'hdb : _GEN_687; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_689 = 8'ha0 == _T_528 ? 8'he0 : _GEN_688; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_690 = 8'ha1 == _T_528 ? 8'h32 : _GEN_689; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_691 = 8'ha2 == _T_528 ? 8'h3a : _GEN_690; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_692 = 8'ha3 == _T_528 ? 8'ha : _GEN_691; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_693 = 8'ha4 == _T_528 ? 8'h49 : _GEN_692; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_694 = 8'ha5 == _T_528 ? 8'h6 : _GEN_693; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_695 = 8'ha6 == _T_528 ? 8'h24 : _GEN_694; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_696 = 8'ha7 == _T_528 ? 8'h5c : _GEN_695; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_697 = 8'ha8 == _T_528 ? 8'hc2 : _GEN_696; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_698 = 8'ha9 == _T_528 ? 8'hd3 : _GEN_697; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_699 = 8'haa == _T_528 ? 8'hac : _GEN_698; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_700 = 8'hab == _T_528 ? 8'h62 : _GEN_699; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_701 = 8'hac == _T_528 ? 8'h91 : _GEN_700; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_702 = 8'had == _T_528 ? 8'h95 : _GEN_701; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_703 = 8'hae == _T_528 ? 8'he4 : _GEN_702; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_704 = 8'haf == _T_528 ? 8'h79 : _GEN_703; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_705 = 8'hb0 == _T_528 ? 8'he7 : _GEN_704; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_706 = 8'hb1 == _T_528 ? 8'hc8 : _GEN_705; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_707 = 8'hb2 == _T_528 ? 8'h37 : _GEN_706; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_708 = 8'hb3 == _T_528 ? 8'h6d : _GEN_707; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_709 = 8'hb4 == _T_528 ? 8'h8d : _GEN_708; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_710 = 8'hb5 == _T_528 ? 8'hd5 : _GEN_709; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_711 = 8'hb6 == _T_528 ? 8'h4e : _GEN_710; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_712 = 8'hb7 == _T_528 ? 8'ha9 : _GEN_711; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_713 = 8'hb8 == _T_528 ? 8'h6c : _GEN_712; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_714 = 8'hb9 == _T_528 ? 8'h56 : _GEN_713; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_715 = 8'hba == _T_528 ? 8'hf4 : _GEN_714; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_716 = 8'hbb == _T_528 ? 8'hea : _GEN_715; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_717 = 8'hbc == _T_528 ? 8'h65 : _GEN_716; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_718 = 8'hbd == _T_528 ? 8'h7a : _GEN_717; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_719 = 8'hbe == _T_528 ? 8'hae : _GEN_718; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_720 = 8'hbf == _T_528 ? 8'h8 : _GEN_719; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_721 = 8'hc0 == _T_528 ? 8'hba : _GEN_720; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_722 = 8'hc1 == _T_528 ? 8'h78 : _GEN_721; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_723 = 8'hc2 == _T_528 ? 8'h25 : _GEN_722; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_724 = 8'hc3 == _T_528 ? 8'h2e : _GEN_723; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_725 = 8'hc4 == _T_528 ? 8'h1c : _GEN_724; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_726 = 8'hc5 == _T_528 ? 8'ha6 : _GEN_725; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_727 = 8'hc6 == _T_528 ? 8'hb4 : _GEN_726; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_728 = 8'hc7 == _T_528 ? 8'hc6 : _GEN_727; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_729 = 8'hc8 == _T_528 ? 8'he8 : _GEN_728; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_730 = 8'hc9 == _T_528 ? 8'hdd : _GEN_729; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_731 = 8'hca == _T_528 ? 8'h74 : _GEN_730; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_732 = 8'hcb == _T_528 ? 8'h1f : _GEN_731; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_733 = 8'hcc == _T_528 ? 8'h4b : _GEN_732; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_734 = 8'hcd == _T_528 ? 8'hbd : _GEN_733; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_735 = 8'hce == _T_528 ? 8'h8b : _GEN_734; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_736 = 8'hcf == _T_528 ? 8'h8a : _GEN_735; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_737 = 8'hd0 == _T_528 ? 8'h70 : _GEN_736; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_738 = 8'hd1 == _T_528 ? 8'h3e : _GEN_737; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_739 = 8'hd2 == _T_528 ? 8'hb5 : _GEN_738; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_740 = 8'hd3 == _T_528 ? 8'h66 : _GEN_739; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_741 = 8'hd4 == _T_528 ? 8'h48 : _GEN_740; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_742 = 8'hd5 == _T_528 ? 8'h3 : _GEN_741; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_743 = 8'hd6 == _T_528 ? 8'hf6 : _GEN_742; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_744 = 8'hd7 == _T_528 ? 8'he : _GEN_743; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_745 = 8'hd8 == _T_528 ? 8'h61 : _GEN_744; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_746 = 8'hd9 == _T_528 ? 8'h35 : _GEN_745; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_747 = 8'hda == _T_528 ? 8'h57 : _GEN_746; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_748 = 8'hdb == _T_528 ? 8'hb9 : _GEN_747; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_749 = 8'hdc == _T_528 ? 8'h86 : _GEN_748; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_750 = 8'hdd == _T_528 ? 8'hc1 : _GEN_749; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_751 = 8'hde == _T_528 ? 8'h1d : _GEN_750; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_752 = 8'hdf == _T_528 ? 8'h9e : _GEN_751; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_753 = 8'he0 == _T_528 ? 8'he1 : _GEN_752; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_754 = 8'he1 == _T_528 ? 8'hf8 : _GEN_753; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_755 = 8'he2 == _T_528 ? 8'h98 : _GEN_754; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_756 = 8'he3 == _T_528 ? 8'h11 : _GEN_755; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_757 = 8'he4 == _T_528 ? 8'h69 : _GEN_756; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_758 = 8'he5 == _T_528 ? 8'hd9 : _GEN_757; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_759 = 8'he6 == _T_528 ? 8'h8e : _GEN_758; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_760 = 8'he7 == _T_528 ? 8'h94 : _GEN_759; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_761 = 8'he8 == _T_528 ? 8'h9b : _GEN_760; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_762 = 8'he9 == _T_528 ? 8'h1e : _GEN_761; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_763 = 8'hea == _T_528 ? 8'h87 : _GEN_762; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_764 = 8'heb == _T_528 ? 8'he9 : _GEN_763; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_765 = 8'hec == _T_528 ? 8'hce : _GEN_764; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_766 = 8'hed == _T_528 ? 8'h55 : _GEN_765; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_767 = 8'hee == _T_528 ? 8'h28 : _GEN_766; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_768 = 8'hef == _T_528 ? 8'hdf : _GEN_767; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_769 = 8'hf0 == _T_528 ? 8'h8c : _GEN_768; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_770 = 8'hf1 == _T_528 ? 8'ha1 : _GEN_769; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_771 = 8'hf2 == _T_528 ? 8'h89 : _GEN_770; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_772 = 8'hf3 == _T_528 ? 8'hd : _GEN_771; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_773 = 8'hf4 == _T_528 ? 8'hbf : _GEN_772; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_774 = 8'hf5 == _T_528 ? 8'he6 : _GEN_773; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_775 = 8'hf6 == _T_528 ? 8'h42 : _GEN_774; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_776 = 8'hf7 == _T_528 ? 8'h68 : _GEN_775; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_777 = 8'hf8 == _T_528 ? 8'h41 : _GEN_776; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_778 = 8'hf9 == _T_528 ? 8'h99 : _GEN_777; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_779 = 8'hfa == _T_528 ? 8'h2d : _GEN_778; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_780 = 8'hfb == _T_528 ? 8'hf : _GEN_779; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_781 = 8'hfc == _T_528 ? 8'hb0 : _GEN_780; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_782 = 8'hfd == _T_528 ? 8'h54 : _GEN_781; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_783 = 8'hfe == _T_528 ? 8'hbb : _GEN_782; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_784 = 8'hff == _T_528 ? 8'h16 : _GEN_783; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_785 = 8'h1 == _T_526 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_786 = 8'h2 == _T_526 ? 8'h77 : _GEN_785; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_787 = 8'h3 == _T_526 ? 8'h7b : _GEN_786; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_788 = 8'h4 == _T_526 ? 8'hf2 : _GEN_787; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_789 = 8'h5 == _T_526 ? 8'h6b : _GEN_788; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_790 = 8'h6 == _T_526 ? 8'h6f : _GEN_789; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_791 = 8'h7 == _T_526 ? 8'hc5 : _GEN_790; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_792 = 8'h8 == _T_526 ? 8'h30 : _GEN_791; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_793 = 8'h9 == _T_526 ? 8'h1 : _GEN_792; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_794 = 8'ha == _T_526 ? 8'h67 : _GEN_793; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_795 = 8'hb == _T_526 ? 8'h2b : _GEN_794; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_796 = 8'hc == _T_526 ? 8'hfe : _GEN_795; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_797 = 8'hd == _T_526 ? 8'hd7 : _GEN_796; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_798 = 8'he == _T_526 ? 8'hab : _GEN_797; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_799 = 8'hf == _T_526 ? 8'h76 : _GEN_798; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_800 = 8'h10 == _T_526 ? 8'hca : _GEN_799; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_801 = 8'h11 == _T_526 ? 8'h82 : _GEN_800; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_802 = 8'h12 == _T_526 ? 8'hc9 : _GEN_801; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_803 = 8'h13 == _T_526 ? 8'h7d : _GEN_802; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_804 = 8'h14 == _T_526 ? 8'hfa : _GEN_803; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_805 = 8'h15 == _T_526 ? 8'h59 : _GEN_804; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_806 = 8'h16 == _T_526 ? 8'h47 : _GEN_805; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_807 = 8'h17 == _T_526 ? 8'hf0 : _GEN_806; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_808 = 8'h18 == _T_526 ? 8'had : _GEN_807; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_809 = 8'h19 == _T_526 ? 8'hd4 : _GEN_808; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_810 = 8'h1a == _T_526 ? 8'ha2 : _GEN_809; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_811 = 8'h1b == _T_526 ? 8'haf : _GEN_810; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_812 = 8'h1c == _T_526 ? 8'h9c : _GEN_811; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_813 = 8'h1d == _T_526 ? 8'ha4 : _GEN_812; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_814 = 8'h1e == _T_526 ? 8'h72 : _GEN_813; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_815 = 8'h1f == _T_526 ? 8'hc0 : _GEN_814; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_816 = 8'h20 == _T_526 ? 8'hb7 : _GEN_815; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_817 = 8'h21 == _T_526 ? 8'hfd : _GEN_816; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_818 = 8'h22 == _T_526 ? 8'h93 : _GEN_817; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_819 = 8'h23 == _T_526 ? 8'h26 : _GEN_818; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_820 = 8'h24 == _T_526 ? 8'h36 : _GEN_819; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_821 = 8'h25 == _T_526 ? 8'h3f : _GEN_820; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_822 = 8'h26 == _T_526 ? 8'hf7 : _GEN_821; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_823 = 8'h27 == _T_526 ? 8'hcc : _GEN_822; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_824 = 8'h28 == _T_526 ? 8'h34 : _GEN_823; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_825 = 8'h29 == _T_526 ? 8'ha5 : _GEN_824; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_826 = 8'h2a == _T_526 ? 8'he5 : _GEN_825; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_827 = 8'h2b == _T_526 ? 8'hf1 : _GEN_826; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_828 = 8'h2c == _T_526 ? 8'h71 : _GEN_827; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_829 = 8'h2d == _T_526 ? 8'hd8 : _GEN_828; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_830 = 8'h2e == _T_526 ? 8'h31 : _GEN_829; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_831 = 8'h2f == _T_526 ? 8'h15 : _GEN_830; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_832 = 8'h30 == _T_526 ? 8'h4 : _GEN_831; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_833 = 8'h31 == _T_526 ? 8'hc7 : _GEN_832; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_834 = 8'h32 == _T_526 ? 8'h23 : _GEN_833; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_835 = 8'h33 == _T_526 ? 8'hc3 : _GEN_834; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_836 = 8'h34 == _T_526 ? 8'h18 : _GEN_835; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_837 = 8'h35 == _T_526 ? 8'h96 : _GEN_836; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_838 = 8'h36 == _T_526 ? 8'h5 : _GEN_837; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_839 = 8'h37 == _T_526 ? 8'h9a : _GEN_838; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_840 = 8'h38 == _T_526 ? 8'h7 : _GEN_839; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_841 = 8'h39 == _T_526 ? 8'h12 : _GEN_840; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_842 = 8'h3a == _T_526 ? 8'h80 : _GEN_841; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_843 = 8'h3b == _T_526 ? 8'he2 : _GEN_842; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_844 = 8'h3c == _T_526 ? 8'heb : _GEN_843; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_845 = 8'h3d == _T_526 ? 8'h27 : _GEN_844; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_846 = 8'h3e == _T_526 ? 8'hb2 : _GEN_845; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_847 = 8'h3f == _T_526 ? 8'h75 : _GEN_846; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_848 = 8'h40 == _T_526 ? 8'h9 : _GEN_847; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_849 = 8'h41 == _T_526 ? 8'h83 : _GEN_848; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_850 = 8'h42 == _T_526 ? 8'h2c : _GEN_849; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_851 = 8'h43 == _T_526 ? 8'h1a : _GEN_850; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_852 = 8'h44 == _T_526 ? 8'h1b : _GEN_851; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_853 = 8'h45 == _T_526 ? 8'h6e : _GEN_852; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_854 = 8'h46 == _T_526 ? 8'h5a : _GEN_853; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_855 = 8'h47 == _T_526 ? 8'ha0 : _GEN_854; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_856 = 8'h48 == _T_526 ? 8'h52 : _GEN_855; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_857 = 8'h49 == _T_526 ? 8'h3b : _GEN_856; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_858 = 8'h4a == _T_526 ? 8'hd6 : _GEN_857; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_859 = 8'h4b == _T_526 ? 8'hb3 : _GEN_858; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_860 = 8'h4c == _T_526 ? 8'h29 : _GEN_859; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_861 = 8'h4d == _T_526 ? 8'he3 : _GEN_860; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_862 = 8'h4e == _T_526 ? 8'h2f : _GEN_861; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_863 = 8'h4f == _T_526 ? 8'h84 : _GEN_862; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_864 = 8'h50 == _T_526 ? 8'h53 : _GEN_863; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_865 = 8'h51 == _T_526 ? 8'hd1 : _GEN_864; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_866 = 8'h52 == _T_526 ? 8'h0 : _GEN_865; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_867 = 8'h53 == _T_526 ? 8'hed : _GEN_866; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_868 = 8'h54 == _T_526 ? 8'h20 : _GEN_867; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_869 = 8'h55 == _T_526 ? 8'hfc : _GEN_868; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_870 = 8'h56 == _T_526 ? 8'hb1 : _GEN_869; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_871 = 8'h57 == _T_526 ? 8'h5b : _GEN_870; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_872 = 8'h58 == _T_526 ? 8'h6a : _GEN_871; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_873 = 8'h59 == _T_526 ? 8'hcb : _GEN_872; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_874 = 8'h5a == _T_526 ? 8'hbe : _GEN_873; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_875 = 8'h5b == _T_526 ? 8'h39 : _GEN_874; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_876 = 8'h5c == _T_526 ? 8'h4a : _GEN_875; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_877 = 8'h5d == _T_526 ? 8'h4c : _GEN_876; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_878 = 8'h5e == _T_526 ? 8'h58 : _GEN_877; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_879 = 8'h5f == _T_526 ? 8'hcf : _GEN_878; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_880 = 8'h60 == _T_526 ? 8'hd0 : _GEN_879; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_881 = 8'h61 == _T_526 ? 8'hef : _GEN_880; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_882 = 8'h62 == _T_526 ? 8'haa : _GEN_881; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_883 = 8'h63 == _T_526 ? 8'hfb : _GEN_882; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_884 = 8'h64 == _T_526 ? 8'h43 : _GEN_883; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_885 = 8'h65 == _T_526 ? 8'h4d : _GEN_884; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_886 = 8'h66 == _T_526 ? 8'h33 : _GEN_885; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_887 = 8'h67 == _T_526 ? 8'h85 : _GEN_886; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_888 = 8'h68 == _T_526 ? 8'h45 : _GEN_887; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_889 = 8'h69 == _T_526 ? 8'hf9 : _GEN_888; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_890 = 8'h6a == _T_526 ? 8'h2 : _GEN_889; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_891 = 8'h6b == _T_526 ? 8'h7f : _GEN_890; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_892 = 8'h6c == _T_526 ? 8'h50 : _GEN_891; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_893 = 8'h6d == _T_526 ? 8'h3c : _GEN_892; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_894 = 8'h6e == _T_526 ? 8'h9f : _GEN_893; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_895 = 8'h6f == _T_526 ? 8'ha8 : _GEN_894; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_896 = 8'h70 == _T_526 ? 8'h51 : _GEN_895; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_897 = 8'h71 == _T_526 ? 8'ha3 : _GEN_896; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_898 = 8'h72 == _T_526 ? 8'h40 : _GEN_897; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_899 = 8'h73 == _T_526 ? 8'h8f : _GEN_898; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_900 = 8'h74 == _T_526 ? 8'h92 : _GEN_899; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_901 = 8'h75 == _T_526 ? 8'h9d : _GEN_900; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_902 = 8'h76 == _T_526 ? 8'h38 : _GEN_901; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_903 = 8'h77 == _T_526 ? 8'hf5 : _GEN_902; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_904 = 8'h78 == _T_526 ? 8'hbc : _GEN_903; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_905 = 8'h79 == _T_526 ? 8'hb6 : _GEN_904; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_906 = 8'h7a == _T_526 ? 8'hda : _GEN_905; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_907 = 8'h7b == _T_526 ? 8'h21 : _GEN_906; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_908 = 8'h7c == _T_526 ? 8'h10 : _GEN_907; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_909 = 8'h7d == _T_526 ? 8'hff : _GEN_908; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_910 = 8'h7e == _T_526 ? 8'hf3 : _GEN_909; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_911 = 8'h7f == _T_526 ? 8'hd2 : _GEN_910; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_912 = 8'h80 == _T_526 ? 8'hcd : _GEN_911; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_913 = 8'h81 == _T_526 ? 8'hc : _GEN_912; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_914 = 8'h82 == _T_526 ? 8'h13 : _GEN_913; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_915 = 8'h83 == _T_526 ? 8'hec : _GEN_914; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_916 = 8'h84 == _T_526 ? 8'h5f : _GEN_915; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_917 = 8'h85 == _T_526 ? 8'h97 : _GEN_916; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_918 = 8'h86 == _T_526 ? 8'h44 : _GEN_917; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_919 = 8'h87 == _T_526 ? 8'h17 : _GEN_918; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_920 = 8'h88 == _T_526 ? 8'hc4 : _GEN_919; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_921 = 8'h89 == _T_526 ? 8'ha7 : _GEN_920; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_922 = 8'h8a == _T_526 ? 8'h7e : _GEN_921; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_923 = 8'h8b == _T_526 ? 8'h3d : _GEN_922; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_924 = 8'h8c == _T_526 ? 8'h64 : _GEN_923; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_925 = 8'h8d == _T_526 ? 8'h5d : _GEN_924; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_926 = 8'h8e == _T_526 ? 8'h19 : _GEN_925; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_927 = 8'h8f == _T_526 ? 8'h73 : _GEN_926; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_928 = 8'h90 == _T_526 ? 8'h60 : _GEN_927; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_929 = 8'h91 == _T_526 ? 8'h81 : _GEN_928; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_930 = 8'h92 == _T_526 ? 8'h4f : _GEN_929; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_931 = 8'h93 == _T_526 ? 8'hdc : _GEN_930; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_932 = 8'h94 == _T_526 ? 8'h22 : _GEN_931; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_933 = 8'h95 == _T_526 ? 8'h2a : _GEN_932; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_934 = 8'h96 == _T_526 ? 8'h90 : _GEN_933; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_935 = 8'h97 == _T_526 ? 8'h88 : _GEN_934; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_936 = 8'h98 == _T_526 ? 8'h46 : _GEN_935; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_937 = 8'h99 == _T_526 ? 8'hee : _GEN_936; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_938 = 8'h9a == _T_526 ? 8'hb8 : _GEN_937; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_939 = 8'h9b == _T_526 ? 8'h14 : _GEN_938; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_940 = 8'h9c == _T_526 ? 8'hde : _GEN_939; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_941 = 8'h9d == _T_526 ? 8'h5e : _GEN_940; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_942 = 8'h9e == _T_526 ? 8'hb : _GEN_941; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_943 = 8'h9f == _T_526 ? 8'hdb : _GEN_942; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_944 = 8'ha0 == _T_526 ? 8'he0 : _GEN_943; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_945 = 8'ha1 == _T_526 ? 8'h32 : _GEN_944; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_946 = 8'ha2 == _T_526 ? 8'h3a : _GEN_945; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_947 = 8'ha3 == _T_526 ? 8'ha : _GEN_946; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_948 = 8'ha4 == _T_526 ? 8'h49 : _GEN_947; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_949 = 8'ha5 == _T_526 ? 8'h6 : _GEN_948; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_950 = 8'ha6 == _T_526 ? 8'h24 : _GEN_949; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_951 = 8'ha7 == _T_526 ? 8'h5c : _GEN_950; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_952 = 8'ha8 == _T_526 ? 8'hc2 : _GEN_951; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_953 = 8'ha9 == _T_526 ? 8'hd3 : _GEN_952; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_954 = 8'haa == _T_526 ? 8'hac : _GEN_953; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_955 = 8'hab == _T_526 ? 8'h62 : _GEN_954; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_956 = 8'hac == _T_526 ? 8'h91 : _GEN_955; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_957 = 8'had == _T_526 ? 8'h95 : _GEN_956; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_958 = 8'hae == _T_526 ? 8'he4 : _GEN_957; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_959 = 8'haf == _T_526 ? 8'h79 : _GEN_958; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_960 = 8'hb0 == _T_526 ? 8'he7 : _GEN_959; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_961 = 8'hb1 == _T_526 ? 8'hc8 : _GEN_960; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_962 = 8'hb2 == _T_526 ? 8'h37 : _GEN_961; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_963 = 8'hb3 == _T_526 ? 8'h6d : _GEN_962; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_964 = 8'hb4 == _T_526 ? 8'h8d : _GEN_963; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_965 = 8'hb5 == _T_526 ? 8'hd5 : _GEN_964; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_966 = 8'hb6 == _T_526 ? 8'h4e : _GEN_965; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_967 = 8'hb7 == _T_526 ? 8'ha9 : _GEN_966; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_968 = 8'hb8 == _T_526 ? 8'h6c : _GEN_967; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_969 = 8'hb9 == _T_526 ? 8'h56 : _GEN_968; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_970 = 8'hba == _T_526 ? 8'hf4 : _GEN_969; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_971 = 8'hbb == _T_526 ? 8'hea : _GEN_970; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_972 = 8'hbc == _T_526 ? 8'h65 : _GEN_971; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_973 = 8'hbd == _T_526 ? 8'h7a : _GEN_972; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_974 = 8'hbe == _T_526 ? 8'hae : _GEN_973; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_975 = 8'hbf == _T_526 ? 8'h8 : _GEN_974; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_976 = 8'hc0 == _T_526 ? 8'hba : _GEN_975; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_977 = 8'hc1 == _T_526 ? 8'h78 : _GEN_976; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_978 = 8'hc2 == _T_526 ? 8'h25 : _GEN_977; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_979 = 8'hc3 == _T_526 ? 8'h2e : _GEN_978; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_980 = 8'hc4 == _T_526 ? 8'h1c : _GEN_979; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_981 = 8'hc5 == _T_526 ? 8'ha6 : _GEN_980; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_982 = 8'hc6 == _T_526 ? 8'hb4 : _GEN_981; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_983 = 8'hc7 == _T_526 ? 8'hc6 : _GEN_982; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_984 = 8'hc8 == _T_526 ? 8'he8 : _GEN_983; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_985 = 8'hc9 == _T_526 ? 8'hdd : _GEN_984; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_986 = 8'hca == _T_526 ? 8'h74 : _GEN_985; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_987 = 8'hcb == _T_526 ? 8'h1f : _GEN_986; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_988 = 8'hcc == _T_526 ? 8'h4b : _GEN_987; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_989 = 8'hcd == _T_526 ? 8'hbd : _GEN_988; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_990 = 8'hce == _T_526 ? 8'h8b : _GEN_989; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_991 = 8'hcf == _T_526 ? 8'h8a : _GEN_990; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_992 = 8'hd0 == _T_526 ? 8'h70 : _GEN_991; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_993 = 8'hd1 == _T_526 ? 8'h3e : _GEN_992; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_994 = 8'hd2 == _T_526 ? 8'hb5 : _GEN_993; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_995 = 8'hd3 == _T_526 ? 8'h66 : _GEN_994; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_996 = 8'hd4 == _T_526 ? 8'h48 : _GEN_995; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_997 = 8'hd5 == _T_526 ? 8'h3 : _GEN_996; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_998 = 8'hd6 == _T_526 ? 8'hf6 : _GEN_997; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_999 = 8'hd7 == _T_526 ? 8'he : _GEN_998; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1000 = 8'hd8 == _T_526 ? 8'h61 : _GEN_999; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1001 = 8'hd9 == _T_526 ? 8'h35 : _GEN_1000; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1002 = 8'hda == _T_526 ? 8'h57 : _GEN_1001; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1003 = 8'hdb == _T_526 ? 8'hb9 : _GEN_1002; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1004 = 8'hdc == _T_526 ? 8'h86 : _GEN_1003; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1005 = 8'hdd == _T_526 ? 8'hc1 : _GEN_1004; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1006 = 8'hde == _T_526 ? 8'h1d : _GEN_1005; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1007 = 8'hdf == _T_526 ? 8'h9e : _GEN_1006; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1008 = 8'he0 == _T_526 ? 8'he1 : _GEN_1007; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1009 = 8'he1 == _T_526 ? 8'hf8 : _GEN_1008; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1010 = 8'he2 == _T_526 ? 8'h98 : _GEN_1009; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1011 = 8'he3 == _T_526 ? 8'h11 : _GEN_1010; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1012 = 8'he4 == _T_526 ? 8'h69 : _GEN_1011; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1013 = 8'he5 == _T_526 ? 8'hd9 : _GEN_1012; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1014 = 8'he6 == _T_526 ? 8'h8e : _GEN_1013; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1015 = 8'he7 == _T_526 ? 8'h94 : _GEN_1014; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1016 = 8'he8 == _T_526 ? 8'h9b : _GEN_1015; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1017 = 8'he9 == _T_526 ? 8'h1e : _GEN_1016; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1018 = 8'hea == _T_526 ? 8'h87 : _GEN_1017; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1019 = 8'heb == _T_526 ? 8'he9 : _GEN_1018; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1020 = 8'hec == _T_526 ? 8'hce : _GEN_1019; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1021 = 8'hed == _T_526 ? 8'h55 : _GEN_1020; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1022 = 8'hee == _T_526 ? 8'h28 : _GEN_1021; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1023 = 8'hef == _T_526 ? 8'hdf : _GEN_1022; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1024 = 8'hf0 == _T_526 ? 8'h8c : _GEN_1023; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1025 = 8'hf1 == _T_526 ? 8'ha1 : _GEN_1024; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1026 = 8'hf2 == _T_526 ? 8'h89 : _GEN_1025; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1027 = 8'hf3 == _T_526 ? 8'hd : _GEN_1026; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1028 = 8'hf4 == _T_526 ? 8'hbf : _GEN_1027; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1029 = 8'hf5 == _T_526 ? 8'he6 : _GEN_1028; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1030 = 8'hf6 == _T_526 ? 8'h42 : _GEN_1029; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1031 = 8'hf7 == _T_526 ? 8'h68 : _GEN_1030; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1032 = 8'hf8 == _T_526 ? 8'h41 : _GEN_1031; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1033 = 8'hf9 == _T_526 ? 8'h99 : _GEN_1032; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1034 = 8'hfa == _T_526 ? 8'h2d : _GEN_1033; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1035 = 8'hfb == _T_526 ? 8'hf : _GEN_1034; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1036 = 8'hfc == _T_526 ? 8'hb0 : _GEN_1035; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1037 = 8'hfd == _T_526 ? 8'h54 : _GEN_1036; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1038 = 8'hfe == _T_526 ? 8'hbb : _GEN_1037; // @[Cat.scala 30:58:@2066.4]
  assign _GEN_1039 = 8'hff == _T_526 ? 8'h16 : _GEN_1038; // @[Cat.scala 30:58:@2066.4]
  assign _T_531 = {_GEN_784,_GEN_1039}; // @[Cat.scala 30:58:@2066.4]
  assign _T_532 = {_T_531,_T_530}; // @[Cat.scala 30:58:@2067.4]
  assign _T_533 = io_addr2[7:0]; // @[sbox.scala 55:25:@2069.4]
  assign _T_535 = io_addr2[15:8]; // @[sbox.scala 56:25:@2070.4]
  assign _T_537 = io_addr2[23:16]; // @[sbox.scala 57:25:@2071.4]
  assign _T_539 = io_addr2[31:24]; // @[sbox.scala 58:25:@2072.4]
  assign _GEN_1040 = 8'h1 == _T_535 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1041 = 8'h2 == _T_535 ? 8'h77 : _GEN_1040; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1042 = 8'h3 == _T_535 ? 8'h7b : _GEN_1041; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1043 = 8'h4 == _T_535 ? 8'hf2 : _GEN_1042; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1044 = 8'h5 == _T_535 ? 8'h6b : _GEN_1043; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1045 = 8'h6 == _T_535 ? 8'h6f : _GEN_1044; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1046 = 8'h7 == _T_535 ? 8'hc5 : _GEN_1045; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1047 = 8'h8 == _T_535 ? 8'h30 : _GEN_1046; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1048 = 8'h9 == _T_535 ? 8'h1 : _GEN_1047; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1049 = 8'ha == _T_535 ? 8'h67 : _GEN_1048; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1050 = 8'hb == _T_535 ? 8'h2b : _GEN_1049; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1051 = 8'hc == _T_535 ? 8'hfe : _GEN_1050; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1052 = 8'hd == _T_535 ? 8'hd7 : _GEN_1051; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1053 = 8'he == _T_535 ? 8'hab : _GEN_1052; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1054 = 8'hf == _T_535 ? 8'h76 : _GEN_1053; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1055 = 8'h10 == _T_535 ? 8'hca : _GEN_1054; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1056 = 8'h11 == _T_535 ? 8'h82 : _GEN_1055; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1057 = 8'h12 == _T_535 ? 8'hc9 : _GEN_1056; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1058 = 8'h13 == _T_535 ? 8'h7d : _GEN_1057; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1059 = 8'h14 == _T_535 ? 8'hfa : _GEN_1058; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1060 = 8'h15 == _T_535 ? 8'h59 : _GEN_1059; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1061 = 8'h16 == _T_535 ? 8'h47 : _GEN_1060; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1062 = 8'h17 == _T_535 ? 8'hf0 : _GEN_1061; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1063 = 8'h18 == _T_535 ? 8'had : _GEN_1062; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1064 = 8'h19 == _T_535 ? 8'hd4 : _GEN_1063; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1065 = 8'h1a == _T_535 ? 8'ha2 : _GEN_1064; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1066 = 8'h1b == _T_535 ? 8'haf : _GEN_1065; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1067 = 8'h1c == _T_535 ? 8'h9c : _GEN_1066; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1068 = 8'h1d == _T_535 ? 8'ha4 : _GEN_1067; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1069 = 8'h1e == _T_535 ? 8'h72 : _GEN_1068; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1070 = 8'h1f == _T_535 ? 8'hc0 : _GEN_1069; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1071 = 8'h20 == _T_535 ? 8'hb7 : _GEN_1070; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1072 = 8'h21 == _T_535 ? 8'hfd : _GEN_1071; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1073 = 8'h22 == _T_535 ? 8'h93 : _GEN_1072; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1074 = 8'h23 == _T_535 ? 8'h26 : _GEN_1073; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1075 = 8'h24 == _T_535 ? 8'h36 : _GEN_1074; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1076 = 8'h25 == _T_535 ? 8'h3f : _GEN_1075; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1077 = 8'h26 == _T_535 ? 8'hf7 : _GEN_1076; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1078 = 8'h27 == _T_535 ? 8'hcc : _GEN_1077; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1079 = 8'h28 == _T_535 ? 8'h34 : _GEN_1078; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1080 = 8'h29 == _T_535 ? 8'ha5 : _GEN_1079; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1081 = 8'h2a == _T_535 ? 8'he5 : _GEN_1080; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1082 = 8'h2b == _T_535 ? 8'hf1 : _GEN_1081; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1083 = 8'h2c == _T_535 ? 8'h71 : _GEN_1082; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1084 = 8'h2d == _T_535 ? 8'hd8 : _GEN_1083; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1085 = 8'h2e == _T_535 ? 8'h31 : _GEN_1084; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1086 = 8'h2f == _T_535 ? 8'h15 : _GEN_1085; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1087 = 8'h30 == _T_535 ? 8'h4 : _GEN_1086; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1088 = 8'h31 == _T_535 ? 8'hc7 : _GEN_1087; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1089 = 8'h32 == _T_535 ? 8'h23 : _GEN_1088; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1090 = 8'h33 == _T_535 ? 8'hc3 : _GEN_1089; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1091 = 8'h34 == _T_535 ? 8'h18 : _GEN_1090; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1092 = 8'h35 == _T_535 ? 8'h96 : _GEN_1091; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1093 = 8'h36 == _T_535 ? 8'h5 : _GEN_1092; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1094 = 8'h37 == _T_535 ? 8'h9a : _GEN_1093; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1095 = 8'h38 == _T_535 ? 8'h7 : _GEN_1094; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1096 = 8'h39 == _T_535 ? 8'h12 : _GEN_1095; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1097 = 8'h3a == _T_535 ? 8'h80 : _GEN_1096; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1098 = 8'h3b == _T_535 ? 8'he2 : _GEN_1097; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1099 = 8'h3c == _T_535 ? 8'heb : _GEN_1098; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1100 = 8'h3d == _T_535 ? 8'h27 : _GEN_1099; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1101 = 8'h3e == _T_535 ? 8'hb2 : _GEN_1100; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1102 = 8'h3f == _T_535 ? 8'h75 : _GEN_1101; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1103 = 8'h40 == _T_535 ? 8'h9 : _GEN_1102; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1104 = 8'h41 == _T_535 ? 8'h83 : _GEN_1103; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1105 = 8'h42 == _T_535 ? 8'h2c : _GEN_1104; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1106 = 8'h43 == _T_535 ? 8'h1a : _GEN_1105; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1107 = 8'h44 == _T_535 ? 8'h1b : _GEN_1106; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1108 = 8'h45 == _T_535 ? 8'h6e : _GEN_1107; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1109 = 8'h46 == _T_535 ? 8'h5a : _GEN_1108; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1110 = 8'h47 == _T_535 ? 8'ha0 : _GEN_1109; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1111 = 8'h48 == _T_535 ? 8'h52 : _GEN_1110; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1112 = 8'h49 == _T_535 ? 8'h3b : _GEN_1111; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1113 = 8'h4a == _T_535 ? 8'hd6 : _GEN_1112; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1114 = 8'h4b == _T_535 ? 8'hb3 : _GEN_1113; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1115 = 8'h4c == _T_535 ? 8'h29 : _GEN_1114; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1116 = 8'h4d == _T_535 ? 8'he3 : _GEN_1115; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1117 = 8'h4e == _T_535 ? 8'h2f : _GEN_1116; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1118 = 8'h4f == _T_535 ? 8'h84 : _GEN_1117; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1119 = 8'h50 == _T_535 ? 8'h53 : _GEN_1118; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1120 = 8'h51 == _T_535 ? 8'hd1 : _GEN_1119; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1121 = 8'h52 == _T_535 ? 8'h0 : _GEN_1120; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1122 = 8'h53 == _T_535 ? 8'hed : _GEN_1121; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1123 = 8'h54 == _T_535 ? 8'h20 : _GEN_1122; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1124 = 8'h55 == _T_535 ? 8'hfc : _GEN_1123; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1125 = 8'h56 == _T_535 ? 8'hb1 : _GEN_1124; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1126 = 8'h57 == _T_535 ? 8'h5b : _GEN_1125; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1127 = 8'h58 == _T_535 ? 8'h6a : _GEN_1126; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1128 = 8'h59 == _T_535 ? 8'hcb : _GEN_1127; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1129 = 8'h5a == _T_535 ? 8'hbe : _GEN_1128; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1130 = 8'h5b == _T_535 ? 8'h39 : _GEN_1129; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1131 = 8'h5c == _T_535 ? 8'h4a : _GEN_1130; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1132 = 8'h5d == _T_535 ? 8'h4c : _GEN_1131; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1133 = 8'h5e == _T_535 ? 8'h58 : _GEN_1132; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1134 = 8'h5f == _T_535 ? 8'hcf : _GEN_1133; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1135 = 8'h60 == _T_535 ? 8'hd0 : _GEN_1134; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1136 = 8'h61 == _T_535 ? 8'hef : _GEN_1135; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1137 = 8'h62 == _T_535 ? 8'haa : _GEN_1136; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1138 = 8'h63 == _T_535 ? 8'hfb : _GEN_1137; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1139 = 8'h64 == _T_535 ? 8'h43 : _GEN_1138; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1140 = 8'h65 == _T_535 ? 8'h4d : _GEN_1139; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1141 = 8'h66 == _T_535 ? 8'h33 : _GEN_1140; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1142 = 8'h67 == _T_535 ? 8'h85 : _GEN_1141; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1143 = 8'h68 == _T_535 ? 8'h45 : _GEN_1142; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1144 = 8'h69 == _T_535 ? 8'hf9 : _GEN_1143; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1145 = 8'h6a == _T_535 ? 8'h2 : _GEN_1144; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1146 = 8'h6b == _T_535 ? 8'h7f : _GEN_1145; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1147 = 8'h6c == _T_535 ? 8'h50 : _GEN_1146; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1148 = 8'h6d == _T_535 ? 8'h3c : _GEN_1147; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1149 = 8'h6e == _T_535 ? 8'h9f : _GEN_1148; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1150 = 8'h6f == _T_535 ? 8'ha8 : _GEN_1149; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1151 = 8'h70 == _T_535 ? 8'h51 : _GEN_1150; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1152 = 8'h71 == _T_535 ? 8'ha3 : _GEN_1151; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1153 = 8'h72 == _T_535 ? 8'h40 : _GEN_1152; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1154 = 8'h73 == _T_535 ? 8'h8f : _GEN_1153; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1155 = 8'h74 == _T_535 ? 8'h92 : _GEN_1154; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1156 = 8'h75 == _T_535 ? 8'h9d : _GEN_1155; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1157 = 8'h76 == _T_535 ? 8'h38 : _GEN_1156; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1158 = 8'h77 == _T_535 ? 8'hf5 : _GEN_1157; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1159 = 8'h78 == _T_535 ? 8'hbc : _GEN_1158; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1160 = 8'h79 == _T_535 ? 8'hb6 : _GEN_1159; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1161 = 8'h7a == _T_535 ? 8'hda : _GEN_1160; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1162 = 8'h7b == _T_535 ? 8'h21 : _GEN_1161; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1163 = 8'h7c == _T_535 ? 8'h10 : _GEN_1162; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1164 = 8'h7d == _T_535 ? 8'hff : _GEN_1163; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1165 = 8'h7e == _T_535 ? 8'hf3 : _GEN_1164; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1166 = 8'h7f == _T_535 ? 8'hd2 : _GEN_1165; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1167 = 8'h80 == _T_535 ? 8'hcd : _GEN_1166; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1168 = 8'h81 == _T_535 ? 8'hc : _GEN_1167; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1169 = 8'h82 == _T_535 ? 8'h13 : _GEN_1168; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1170 = 8'h83 == _T_535 ? 8'hec : _GEN_1169; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1171 = 8'h84 == _T_535 ? 8'h5f : _GEN_1170; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1172 = 8'h85 == _T_535 ? 8'h97 : _GEN_1171; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1173 = 8'h86 == _T_535 ? 8'h44 : _GEN_1172; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1174 = 8'h87 == _T_535 ? 8'h17 : _GEN_1173; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1175 = 8'h88 == _T_535 ? 8'hc4 : _GEN_1174; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1176 = 8'h89 == _T_535 ? 8'ha7 : _GEN_1175; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1177 = 8'h8a == _T_535 ? 8'h7e : _GEN_1176; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1178 = 8'h8b == _T_535 ? 8'h3d : _GEN_1177; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1179 = 8'h8c == _T_535 ? 8'h64 : _GEN_1178; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1180 = 8'h8d == _T_535 ? 8'h5d : _GEN_1179; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1181 = 8'h8e == _T_535 ? 8'h19 : _GEN_1180; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1182 = 8'h8f == _T_535 ? 8'h73 : _GEN_1181; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1183 = 8'h90 == _T_535 ? 8'h60 : _GEN_1182; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1184 = 8'h91 == _T_535 ? 8'h81 : _GEN_1183; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1185 = 8'h92 == _T_535 ? 8'h4f : _GEN_1184; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1186 = 8'h93 == _T_535 ? 8'hdc : _GEN_1185; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1187 = 8'h94 == _T_535 ? 8'h22 : _GEN_1186; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1188 = 8'h95 == _T_535 ? 8'h2a : _GEN_1187; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1189 = 8'h96 == _T_535 ? 8'h90 : _GEN_1188; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1190 = 8'h97 == _T_535 ? 8'h88 : _GEN_1189; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1191 = 8'h98 == _T_535 ? 8'h46 : _GEN_1190; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1192 = 8'h99 == _T_535 ? 8'hee : _GEN_1191; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1193 = 8'h9a == _T_535 ? 8'hb8 : _GEN_1192; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1194 = 8'h9b == _T_535 ? 8'h14 : _GEN_1193; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1195 = 8'h9c == _T_535 ? 8'hde : _GEN_1194; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1196 = 8'h9d == _T_535 ? 8'h5e : _GEN_1195; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1197 = 8'h9e == _T_535 ? 8'hb : _GEN_1196; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1198 = 8'h9f == _T_535 ? 8'hdb : _GEN_1197; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1199 = 8'ha0 == _T_535 ? 8'he0 : _GEN_1198; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1200 = 8'ha1 == _T_535 ? 8'h32 : _GEN_1199; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1201 = 8'ha2 == _T_535 ? 8'h3a : _GEN_1200; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1202 = 8'ha3 == _T_535 ? 8'ha : _GEN_1201; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1203 = 8'ha4 == _T_535 ? 8'h49 : _GEN_1202; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1204 = 8'ha5 == _T_535 ? 8'h6 : _GEN_1203; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1205 = 8'ha6 == _T_535 ? 8'h24 : _GEN_1204; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1206 = 8'ha7 == _T_535 ? 8'h5c : _GEN_1205; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1207 = 8'ha8 == _T_535 ? 8'hc2 : _GEN_1206; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1208 = 8'ha9 == _T_535 ? 8'hd3 : _GEN_1207; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1209 = 8'haa == _T_535 ? 8'hac : _GEN_1208; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1210 = 8'hab == _T_535 ? 8'h62 : _GEN_1209; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1211 = 8'hac == _T_535 ? 8'h91 : _GEN_1210; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1212 = 8'had == _T_535 ? 8'h95 : _GEN_1211; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1213 = 8'hae == _T_535 ? 8'he4 : _GEN_1212; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1214 = 8'haf == _T_535 ? 8'h79 : _GEN_1213; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1215 = 8'hb0 == _T_535 ? 8'he7 : _GEN_1214; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1216 = 8'hb1 == _T_535 ? 8'hc8 : _GEN_1215; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1217 = 8'hb2 == _T_535 ? 8'h37 : _GEN_1216; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1218 = 8'hb3 == _T_535 ? 8'h6d : _GEN_1217; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1219 = 8'hb4 == _T_535 ? 8'h8d : _GEN_1218; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1220 = 8'hb5 == _T_535 ? 8'hd5 : _GEN_1219; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1221 = 8'hb6 == _T_535 ? 8'h4e : _GEN_1220; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1222 = 8'hb7 == _T_535 ? 8'ha9 : _GEN_1221; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1223 = 8'hb8 == _T_535 ? 8'h6c : _GEN_1222; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1224 = 8'hb9 == _T_535 ? 8'h56 : _GEN_1223; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1225 = 8'hba == _T_535 ? 8'hf4 : _GEN_1224; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1226 = 8'hbb == _T_535 ? 8'hea : _GEN_1225; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1227 = 8'hbc == _T_535 ? 8'h65 : _GEN_1226; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1228 = 8'hbd == _T_535 ? 8'h7a : _GEN_1227; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1229 = 8'hbe == _T_535 ? 8'hae : _GEN_1228; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1230 = 8'hbf == _T_535 ? 8'h8 : _GEN_1229; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1231 = 8'hc0 == _T_535 ? 8'hba : _GEN_1230; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1232 = 8'hc1 == _T_535 ? 8'h78 : _GEN_1231; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1233 = 8'hc2 == _T_535 ? 8'h25 : _GEN_1232; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1234 = 8'hc3 == _T_535 ? 8'h2e : _GEN_1233; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1235 = 8'hc4 == _T_535 ? 8'h1c : _GEN_1234; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1236 = 8'hc5 == _T_535 ? 8'ha6 : _GEN_1235; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1237 = 8'hc6 == _T_535 ? 8'hb4 : _GEN_1236; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1238 = 8'hc7 == _T_535 ? 8'hc6 : _GEN_1237; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1239 = 8'hc8 == _T_535 ? 8'he8 : _GEN_1238; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1240 = 8'hc9 == _T_535 ? 8'hdd : _GEN_1239; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1241 = 8'hca == _T_535 ? 8'h74 : _GEN_1240; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1242 = 8'hcb == _T_535 ? 8'h1f : _GEN_1241; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1243 = 8'hcc == _T_535 ? 8'h4b : _GEN_1242; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1244 = 8'hcd == _T_535 ? 8'hbd : _GEN_1243; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1245 = 8'hce == _T_535 ? 8'h8b : _GEN_1244; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1246 = 8'hcf == _T_535 ? 8'h8a : _GEN_1245; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1247 = 8'hd0 == _T_535 ? 8'h70 : _GEN_1246; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1248 = 8'hd1 == _T_535 ? 8'h3e : _GEN_1247; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1249 = 8'hd2 == _T_535 ? 8'hb5 : _GEN_1248; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1250 = 8'hd3 == _T_535 ? 8'h66 : _GEN_1249; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1251 = 8'hd4 == _T_535 ? 8'h48 : _GEN_1250; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1252 = 8'hd5 == _T_535 ? 8'h3 : _GEN_1251; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1253 = 8'hd6 == _T_535 ? 8'hf6 : _GEN_1252; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1254 = 8'hd7 == _T_535 ? 8'he : _GEN_1253; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1255 = 8'hd8 == _T_535 ? 8'h61 : _GEN_1254; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1256 = 8'hd9 == _T_535 ? 8'h35 : _GEN_1255; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1257 = 8'hda == _T_535 ? 8'h57 : _GEN_1256; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1258 = 8'hdb == _T_535 ? 8'hb9 : _GEN_1257; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1259 = 8'hdc == _T_535 ? 8'h86 : _GEN_1258; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1260 = 8'hdd == _T_535 ? 8'hc1 : _GEN_1259; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1261 = 8'hde == _T_535 ? 8'h1d : _GEN_1260; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1262 = 8'hdf == _T_535 ? 8'h9e : _GEN_1261; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1263 = 8'he0 == _T_535 ? 8'he1 : _GEN_1262; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1264 = 8'he1 == _T_535 ? 8'hf8 : _GEN_1263; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1265 = 8'he2 == _T_535 ? 8'h98 : _GEN_1264; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1266 = 8'he3 == _T_535 ? 8'h11 : _GEN_1265; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1267 = 8'he4 == _T_535 ? 8'h69 : _GEN_1266; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1268 = 8'he5 == _T_535 ? 8'hd9 : _GEN_1267; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1269 = 8'he6 == _T_535 ? 8'h8e : _GEN_1268; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1270 = 8'he7 == _T_535 ? 8'h94 : _GEN_1269; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1271 = 8'he8 == _T_535 ? 8'h9b : _GEN_1270; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1272 = 8'he9 == _T_535 ? 8'h1e : _GEN_1271; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1273 = 8'hea == _T_535 ? 8'h87 : _GEN_1272; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1274 = 8'heb == _T_535 ? 8'he9 : _GEN_1273; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1275 = 8'hec == _T_535 ? 8'hce : _GEN_1274; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1276 = 8'hed == _T_535 ? 8'h55 : _GEN_1275; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1277 = 8'hee == _T_535 ? 8'h28 : _GEN_1276; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1278 = 8'hef == _T_535 ? 8'hdf : _GEN_1277; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1279 = 8'hf0 == _T_535 ? 8'h8c : _GEN_1278; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1280 = 8'hf1 == _T_535 ? 8'ha1 : _GEN_1279; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1281 = 8'hf2 == _T_535 ? 8'h89 : _GEN_1280; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1282 = 8'hf3 == _T_535 ? 8'hd : _GEN_1281; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1283 = 8'hf4 == _T_535 ? 8'hbf : _GEN_1282; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1284 = 8'hf5 == _T_535 ? 8'he6 : _GEN_1283; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1285 = 8'hf6 == _T_535 ? 8'h42 : _GEN_1284; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1286 = 8'hf7 == _T_535 ? 8'h68 : _GEN_1285; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1287 = 8'hf8 == _T_535 ? 8'h41 : _GEN_1286; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1288 = 8'hf9 == _T_535 ? 8'h99 : _GEN_1287; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1289 = 8'hfa == _T_535 ? 8'h2d : _GEN_1288; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1290 = 8'hfb == _T_535 ? 8'hf : _GEN_1289; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1291 = 8'hfc == _T_535 ? 8'hb0 : _GEN_1290; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1292 = 8'hfd == _T_535 ? 8'h54 : _GEN_1291; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1293 = 8'hfe == _T_535 ? 8'hbb : _GEN_1292; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1294 = 8'hff == _T_535 ? 8'h16 : _GEN_1293; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1295 = 8'h1 == _T_533 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1296 = 8'h2 == _T_533 ? 8'h77 : _GEN_1295; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1297 = 8'h3 == _T_533 ? 8'h7b : _GEN_1296; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1298 = 8'h4 == _T_533 ? 8'hf2 : _GEN_1297; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1299 = 8'h5 == _T_533 ? 8'h6b : _GEN_1298; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1300 = 8'h6 == _T_533 ? 8'h6f : _GEN_1299; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1301 = 8'h7 == _T_533 ? 8'hc5 : _GEN_1300; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1302 = 8'h8 == _T_533 ? 8'h30 : _GEN_1301; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1303 = 8'h9 == _T_533 ? 8'h1 : _GEN_1302; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1304 = 8'ha == _T_533 ? 8'h67 : _GEN_1303; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1305 = 8'hb == _T_533 ? 8'h2b : _GEN_1304; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1306 = 8'hc == _T_533 ? 8'hfe : _GEN_1305; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1307 = 8'hd == _T_533 ? 8'hd7 : _GEN_1306; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1308 = 8'he == _T_533 ? 8'hab : _GEN_1307; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1309 = 8'hf == _T_533 ? 8'h76 : _GEN_1308; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1310 = 8'h10 == _T_533 ? 8'hca : _GEN_1309; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1311 = 8'h11 == _T_533 ? 8'h82 : _GEN_1310; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1312 = 8'h12 == _T_533 ? 8'hc9 : _GEN_1311; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1313 = 8'h13 == _T_533 ? 8'h7d : _GEN_1312; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1314 = 8'h14 == _T_533 ? 8'hfa : _GEN_1313; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1315 = 8'h15 == _T_533 ? 8'h59 : _GEN_1314; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1316 = 8'h16 == _T_533 ? 8'h47 : _GEN_1315; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1317 = 8'h17 == _T_533 ? 8'hf0 : _GEN_1316; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1318 = 8'h18 == _T_533 ? 8'had : _GEN_1317; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1319 = 8'h19 == _T_533 ? 8'hd4 : _GEN_1318; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1320 = 8'h1a == _T_533 ? 8'ha2 : _GEN_1319; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1321 = 8'h1b == _T_533 ? 8'haf : _GEN_1320; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1322 = 8'h1c == _T_533 ? 8'h9c : _GEN_1321; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1323 = 8'h1d == _T_533 ? 8'ha4 : _GEN_1322; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1324 = 8'h1e == _T_533 ? 8'h72 : _GEN_1323; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1325 = 8'h1f == _T_533 ? 8'hc0 : _GEN_1324; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1326 = 8'h20 == _T_533 ? 8'hb7 : _GEN_1325; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1327 = 8'h21 == _T_533 ? 8'hfd : _GEN_1326; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1328 = 8'h22 == _T_533 ? 8'h93 : _GEN_1327; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1329 = 8'h23 == _T_533 ? 8'h26 : _GEN_1328; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1330 = 8'h24 == _T_533 ? 8'h36 : _GEN_1329; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1331 = 8'h25 == _T_533 ? 8'h3f : _GEN_1330; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1332 = 8'h26 == _T_533 ? 8'hf7 : _GEN_1331; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1333 = 8'h27 == _T_533 ? 8'hcc : _GEN_1332; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1334 = 8'h28 == _T_533 ? 8'h34 : _GEN_1333; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1335 = 8'h29 == _T_533 ? 8'ha5 : _GEN_1334; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1336 = 8'h2a == _T_533 ? 8'he5 : _GEN_1335; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1337 = 8'h2b == _T_533 ? 8'hf1 : _GEN_1336; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1338 = 8'h2c == _T_533 ? 8'h71 : _GEN_1337; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1339 = 8'h2d == _T_533 ? 8'hd8 : _GEN_1338; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1340 = 8'h2e == _T_533 ? 8'h31 : _GEN_1339; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1341 = 8'h2f == _T_533 ? 8'h15 : _GEN_1340; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1342 = 8'h30 == _T_533 ? 8'h4 : _GEN_1341; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1343 = 8'h31 == _T_533 ? 8'hc7 : _GEN_1342; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1344 = 8'h32 == _T_533 ? 8'h23 : _GEN_1343; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1345 = 8'h33 == _T_533 ? 8'hc3 : _GEN_1344; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1346 = 8'h34 == _T_533 ? 8'h18 : _GEN_1345; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1347 = 8'h35 == _T_533 ? 8'h96 : _GEN_1346; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1348 = 8'h36 == _T_533 ? 8'h5 : _GEN_1347; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1349 = 8'h37 == _T_533 ? 8'h9a : _GEN_1348; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1350 = 8'h38 == _T_533 ? 8'h7 : _GEN_1349; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1351 = 8'h39 == _T_533 ? 8'h12 : _GEN_1350; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1352 = 8'h3a == _T_533 ? 8'h80 : _GEN_1351; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1353 = 8'h3b == _T_533 ? 8'he2 : _GEN_1352; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1354 = 8'h3c == _T_533 ? 8'heb : _GEN_1353; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1355 = 8'h3d == _T_533 ? 8'h27 : _GEN_1354; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1356 = 8'h3e == _T_533 ? 8'hb2 : _GEN_1355; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1357 = 8'h3f == _T_533 ? 8'h75 : _GEN_1356; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1358 = 8'h40 == _T_533 ? 8'h9 : _GEN_1357; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1359 = 8'h41 == _T_533 ? 8'h83 : _GEN_1358; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1360 = 8'h42 == _T_533 ? 8'h2c : _GEN_1359; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1361 = 8'h43 == _T_533 ? 8'h1a : _GEN_1360; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1362 = 8'h44 == _T_533 ? 8'h1b : _GEN_1361; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1363 = 8'h45 == _T_533 ? 8'h6e : _GEN_1362; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1364 = 8'h46 == _T_533 ? 8'h5a : _GEN_1363; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1365 = 8'h47 == _T_533 ? 8'ha0 : _GEN_1364; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1366 = 8'h48 == _T_533 ? 8'h52 : _GEN_1365; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1367 = 8'h49 == _T_533 ? 8'h3b : _GEN_1366; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1368 = 8'h4a == _T_533 ? 8'hd6 : _GEN_1367; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1369 = 8'h4b == _T_533 ? 8'hb3 : _GEN_1368; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1370 = 8'h4c == _T_533 ? 8'h29 : _GEN_1369; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1371 = 8'h4d == _T_533 ? 8'he3 : _GEN_1370; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1372 = 8'h4e == _T_533 ? 8'h2f : _GEN_1371; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1373 = 8'h4f == _T_533 ? 8'h84 : _GEN_1372; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1374 = 8'h50 == _T_533 ? 8'h53 : _GEN_1373; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1375 = 8'h51 == _T_533 ? 8'hd1 : _GEN_1374; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1376 = 8'h52 == _T_533 ? 8'h0 : _GEN_1375; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1377 = 8'h53 == _T_533 ? 8'hed : _GEN_1376; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1378 = 8'h54 == _T_533 ? 8'h20 : _GEN_1377; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1379 = 8'h55 == _T_533 ? 8'hfc : _GEN_1378; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1380 = 8'h56 == _T_533 ? 8'hb1 : _GEN_1379; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1381 = 8'h57 == _T_533 ? 8'h5b : _GEN_1380; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1382 = 8'h58 == _T_533 ? 8'h6a : _GEN_1381; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1383 = 8'h59 == _T_533 ? 8'hcb : _GEN_1382; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1384 = 8'h5a == _T_533 ? 8'hbe : _GEN_1383; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1385 = 8'h5b == _T_533 ? 8'h39 : _GEN_1384; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1386 = 8'h5c == _T_533 ? 8'h4a : _GEN_1385; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1387 = 8'h5d == _T_533 ? 8'h4c : _GEN_1386; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1388 = 8'h5e == _T_533 ? 8'h58 : _GEN_1387; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1389 = 8'h5f == _T_533 ? 8'hcf : _GEN_1388; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1390 = 8'h60 == _T_533 ? 8'hd0 : _GEN_1389; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1391 = 8'h61 == _T_533 ? 8'hef : _GEN_1390; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1392 = 8'h62 == _T_533 ? 8'haa : _GEN_1391; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1393 = 8'h63 == _T_533 ? 8'hfb : _GEN_1392; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1394 = 8'h64 == _T_533 ? 8'h43 : _GEN_1393; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1395 = 8'h65 == _T_533 ? 8'h4d : _GEN_1394; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1396 = 8'h66 == _T_533 ? 8'h33 : _GEN_1395; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1397 = 8'h67 == _T_533 ? 8'h85 : _GEN_1396; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1398 = 8'h68 == _T_533 ? 8'h45 : _GEN_1397; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1399 = 8'h69 == _T_533 ? 8'hf9 : _GEN_1398; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1400 = 8'h6a == _T_533 ? 8'h2 : _GEN_1399; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1401 = 8'h6b == _T_533 ? 8'h7f : _GEN_1400; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1402 = 8'h6c == _T_533 ? 8'h50 : _GEN_1401; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1403 = 8'h6d == _T_533 ? 8'h3c : _GEN_1402; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1404 = 8'h6e == _T_533 ? 8'h9f : _GEN_1403; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1405 = 8'h6f == _T_533 ? 8'ha8 : _GEN_1404; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1406 = 8'h70 == _T_533 ? 8'h51 : _GEN_1405; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1407 = 8'h71 == _T_533 ? 8'ha3 : _GEN_1406; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1408 = 8'h72 == _T_533 ? 8'h40 : _GEN_1407; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1409 = 8'h73 == _T_533 ? 8'h8f : _GEN_1408; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1410 = 8'h74 == _T_533 ? 8'h92 : _GEN_1409; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1411 = 8'h75 == _T_533 ? 8'h9d : _GEN_1410; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1412 = 8'h76 == _T_533 ? 8'h38 : _GEN_1411; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1413 = 8'h77 == _T_533 ? 8'hf5 : _GEN_1412; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1414 = 8'h78 == _T_533 ? 8'hbc : _GEN_1413; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1415 = 8'h79 == _T_533 ? 8'hb6 : _GEN_1414; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1416 = 8'h7a == _T_533 ? 8'hda : _GEN_1415; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1417 = 8'h7b == _T_533 ? 8'h21 : _GEN_1416; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1418 = 8'h7c == _T_533 ? 8'h10 : _GEN_1417; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1419 = 8'h7d == _T_533 ? 8'hff : _GEN_1418; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1420 = 8'h7e == _T_533 ? 8'hf3 : _GEN_1419; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1421 = 8'h7f == _T_533 ? 8'hd2 : _GEN_1420; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1422 = 8'h80 == _T_533 ? 8'hcd : _GEN_1421; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1423 = 8'h81 == _T_533 ? 8'hc : _GEN_1422; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1424 = 8'h82 == _T_533 ? 8'h13 : _GEN_1423; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1425 = 8'h83 == _T_533 ? 8'hec : _GEN_1424; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1426 = 8'h84 == _T_533 ? 8'h5f : _GEN_1425; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1427 = 8'h85 == _T_533 ? 8'h97 : _GEN_1426; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1428 = 8'h86 == _T_533 ? 8'h44 : _GEN_1427; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1429 = 8'h87 == _T_533 ? 8'h17 : _GEN_1428; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1430 = 8'h88 == _T_533 ? 8'hc4 : _GEN_1429; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1431 = 8'h89 == _T_533 ? 8'ha7 : _GEN_1430; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1432 = 8'h8a == _T_533 ? 8'h7e : _GEN_1431; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1433 = 8'h8b == _T_533 ? 8'h3d : _GEN_1432; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1434 = 8'h8c == _T_533 ? 8'h64 : _GEN_1433; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1435 = 8'h8d == _T_533 ? 8'h5d : _GEN_1434; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1436 = 8'h8e == _T_533 ? 8'h19 : _GEN_1435; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1437 = 8'h8f == _T_533 ? 8'h73 : _GEN_1436; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1438 = 8'h90 == _T_533 ? 8'h60 : _GEN_1437; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1439 = 8'h91 == _T_533 ? 8'h81 : _GEN_1438; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1440 = 8'h92 == _T_533 ? 8'h4f : _GEN_1439; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1441 = 8'h93 == _T_533 ? 8'hdc : _GEN_1440; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1442 = 8'h94 == _T_533 ? 8'h22 : _GEN_1441; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1443 = 8'h95 == _T_533 ? 8'h2a : _GEN_1442; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1444 = 8'h96 == _T_533 ? 8'h90 : _GEN_1443; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1445 = 8'h97 == _T_533 ? 8'h88 : _GEN_1444; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1446 = 8'h98 == _T_533 ? 8'h46 : _GEN_1445; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1447 = 8'h99 == _T_533 ? 8'hee : _GEN_1446; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1448 = 8'h9a == _T_533 ? 8'hb8 : _GEN_1447; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1449 = 8'h9b == _T_533 ? 8'h14 : _GEN_1448; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1450 = 8'h9c == _T_533 ? 8'hde : _GEN_1449; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1451 = 8'h9d == _T_533 ? 8'h5e : _GEN_1450; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1452 = 8'h9e == _T_533 ? 8'hb : _GEN_1451; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1453 = 8'h9f == _T_533 ? 8'hdb : _GEN_1452; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1454 = 8'ha0 == _T_533 ? 8'he0 : _GEN_1453; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1455 = 8'ha1 == _T_533 ? 8'h32 : _GEN_1454; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1456 = 8'ha2 == _T_533 ? 8'h3a : _GEN_1455; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1457 = 8'ha3 == _T_533 ? 8'ha : _GEN_1456; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1458 = 8'ha4 == _T_533 ? 8'h49 : _GEN_1457; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1459 = 8'ha5 == _T_533 ? 8'h6 : _GEN_1458; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1460 = 8'ha6 == _T_533 ? 8'h24 : _GEN_1459; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1461 = 8'ha7 == _T_533 ? 8'h5c : _GEN_1460; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1462 = 8'ha8 == _T_533 ? 8'hc2 : _GEN_1461; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1463 = 8'ha9 == _T_533 ? 8'hd3 : _GEN_1462; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1464 = 8'haa == _T_533 ? 8'hac : _GEN_1463; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1465 = 8'hab == _T_533 ? 8'h62 : _GEN_1464; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1466 = 8'hac == _T_533 ? 8'h91 : _GEN_1465; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1467 = 8'had == _T_533 ? 8'h95 : _GEN_1466; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1468 = 8'hae == _T_533 ? 8'he4 : _GEN_1467; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1469 = 8'haf == _T_533 ? 8'h79 : _GEN_1468; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1470 = 8'hb0 == _T_533 ? 8'he7 : _GEN_1469; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1471 = 8'hb1 == _T_533 ? 8'hc8 : _GEN_1470; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1472 = 8'hb2 == _T_533 ? 8'h37 : _GEN_1471; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1473 = 8'hb3 == _T_533 ? 8'h6d : _GEN_1472; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1474 = 8'hb4 == _T_533 ? 8'h8d : _GEN_1473; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1475 = 8'hb5 == _T_533 ? 8'hd5 : _GEN_1474; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1476 = 8'hb6 == _T_533 ? 8'h4e : _GEN_1475; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1477 = 8'hb7 == _T_533 ? 8'ha9 : _GEN_1476; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1478 = 8'hb8 == _T_533 ? 8'h6c : _GEN_1477; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1479 = 8'hb9 == _T_533 ? 8'h56 : _GEN_1478; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1480 = 8'hba == _T_533 ? 8'hf4 : _GEN_1479; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1481 = 8'hbb == _T_533 ? 8'hea : _GEN_1480; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1482 = 8'hbc == _T_533 ? 8'h65 : _GEN_1481; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1483 = 8'hbd == _T_533 ? 8'h7a : _GEN_1482; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1484 = 8'hbe == _T_533 ? 8'hae : _GEN_1483; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1485 = 8'hbf == _T_533 ? 8'h8 : _GEN_1484; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1486 = 8'hc0 == _T_533 ? 8'hba : _GEN_1485; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1487 = 8'hc1 == _T_533 ? 8'h78 : _GEN_1486; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1488 = 8'hc2 == _T_533 ? 8'h25 : _GEN_1487; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1489 = 8'hc3 == _T_533 ? 8'h2e : _GEN_1488; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1490 = 8'hc4 == _T_533 ? 8'h1c : _GEN_1489; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1491 = 8'hc5 == _T_533 ? 8'ha6 : _GEN_1490; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1492 = 8'hc6 == _T_533 ? 8'hb4 : _GEN_1491; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1493 = 8'hc7 == _T_533 ? 8'hc6 : _GEN_1492; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1494 = 8'hc8 == _T_533 ? 8'he8 : _GEN_1493; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1495 = 8'hc9 == _T_533 ? 8'hdd : _GEN_1494; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1496 = 8'hca == _T_533 ? 8'h74 : _GEN_1495; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1497 = 8'hcb == _T_533 ? 8'h1f : _GEN_1496; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1498 = 8'hcc == _T_533 ? 8'h4b : _GEN_1497; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1499 = 8'hcd == _T_533 ? 8'hbd : _GEN_1498; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1500 = 8'hce == _T_533 ? 8'h8b : _GEN_1499; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1501 = 8'hcf == _T_533 ? 8'h8a : _GEN_1500; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1502 = 8'hd0 == _T_533 ? 8'h70 : _GEN_1501; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1503 = 8'hd1 == _T_533 ? 8'h3e : _GEN_1502; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1504 = 8'hd2 == _T_533 ? 8'hb5 : _GEN_1503; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1505 = 8'hd3 == _T_533 ? 8'h66 : _GEN_1504; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1506 = 8'hd4 == _T_533 ? 8'h48 : _GEN_1505; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1507 = 8'hd5 == _T_533 ? 8'h3 : _GEN_1506; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1508 = 8'hd6 == _T_533 ? 8'hf6 : _GEN_1507; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1509 = 8'hd7 == _T_533 ? 8'he : _GEN_1508; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1510 = 8'hd8 == _T_533 ? 8'h61 : _GEN_1509; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1511 = 8'hd9 == _T_533 ? 8'h35 : _GEN_1510; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1512 = 8'hda == _T_533 ? 8'h57 : _GEN_1511; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1513 = 8'hdb == _T_533 ? 8'hb9 : _GEN_1512; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1514 = 8'hdc == _T_533 ? 8'h86 : _GEN_1513; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1515 = 8'hdd == _T_533 ? 8'hc1 : _GEN_1514; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1516 = 8'hde == _T_533 ? 8'h1d : _GEN_1515; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1517 = 8'hdf == _T_533 ? 8'h9e : _GEN_1516; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1518 = 8'he0 == _T_533 ? 8'he1 : _GEN_1517; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1519 = 8'he1 == _T_533 ? 8'hf8 : _GEN_1518; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1520 = 8'he2 == _T_533 ? 8'h98 : _GEN_1519; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1521 = 8'he3 == _T_533 ? 8'h11 : _GEN_1520; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1522 = 8'he4 == _T_533 ? 8'h69 : _GEN_1521; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1523 = 8'he5 == _T_533 ? 8'hd9 : _GEN_1522; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1524 = 8'he6 == _T_533 ? 8'h8e : _GEN_1523; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1525 = 8'he7 == _T_533 ? 8'h94 : _GEN_1524; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1526 = 8'he8 == _T_533 ? 8'h9b : _GEN_1525; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1527 = 8'he9 == _T_533 ? 8'h1e : _GEN_1526; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1528 = 8'hea == _T_533 ? 8'h87 : _GEN_1527; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1529 = 8'heb == _T_533 ? 8'he9 : _GEN_1528; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1530 = 8'hec == _T_533 ? 8'hce : _GEN_1529; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1531 = 8'hed == _T_533 ? 8'h55 : _GEN_1530; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1532 = 8'hee == _T_533 ? 8'h28 : _GEN_1531; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1533 = 8'hef == _T_533 ? 8'hdf : _GEN_1532; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1534 = 8'hf0 == _T_533 ? 8'h8c : _GEN_1533; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1535 = 8'hf1 == _T_533 ? 8'ha1 : _GEN_1534; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1536 = 8'hf2 == _T_533 ? 8'h89 : _GEN_1535; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1537 = 8'hf3 == _T_533 ? 8'hd : _GEN_1536; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1538 = 8'hf4 == _T_533 ? 8'hbf : _GEN_1537; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1539 = 8'hf5 == _T_533 ? 8'he6 : _GEN_1538; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1540 = 8'hf6 == _T_533 ? 8'h42 : _GEN_1539; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1541 = 8'hf7 == _T_533 ? 8'h68 : _GEN_1540; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1542 = 8'hf8 == _T_533 ? 8'h41 : _GEN_1541; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1543 = 8'hf9 == _T_533 ? 8'h99 : _GEN_1542; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1544 = 8'hfa == _T_533 ? 8'h2d : _GEN_1543; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1545 = 8'hfb == _T_533 ? 8'hf : _GEN_1544; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1546 = 8'hfc == _T_533 ? 8'hb0 : _GEN_1545; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1547 = 8'hfd == _T_533 ? 8'h54 : _GEN_1546; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1548 = 8'hfe == _T_533 ? 8'hbb : _GEN_1547; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1549 = 8'hff == _T_533 ? 8'h16 : _GEN_1548; // @[Cat.scala 30:58:@2073.4]
  assign _T_541 = {_GEN_1294,_GEN_1549}; // @[Cat.scala 30:58:@2073.4]
  assign _GEN_1550 = 8'h1 == _T_539 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1551 = 8'h2 == _T_539 ? 8'h77 : _GEN_1550; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1552 = 8'h3 == _T_539 ? 8'h7b : _GEN_1551; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1553 = 8'h4 == _T_539 ? 8'hf2 : _GEN_1552; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1554 = 8'h5 == _T_539 ? 8'h6b : _GEN_1553; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1555 = 8'h6 == _T_539 ? 8'h6f : _GEN_1554; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1556 = 8'h7 == _T_539 ? 8'hc5 : _GEN_1555; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1557 = 8'h8 == _T_539 ? 8'h30 : _GEN_1556; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1558 = 8'h9 == _T_539 ? 8'h1 : _GEN_1557; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1559 = 8'ha == _T_539 ? 8'h67 : _GEN_1558; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1560 = 8'hb == _T_539 ? 8'h2b : _GEN_1559; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1561 = 8'hc == _T_539 ? 8'hfe : _GEN_1560; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1562 = 8'hd == _T_539 ? 8'hd7 : _GEN_1561; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1563 = 8'he == _T_539 ? 8'hab : _GEN_1562; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1564 = 8'hf == _T_539 ? 8'h76 : _GEN_1563; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1565 = 8'h10 == _T_539 ? 8'hca : _GEN_1564; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1566 = 8'h11 == _T_539 ? 8'h82 : _GEN_1565; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1567 = 8'h12 == _T_539 ? 8'hc9 : _GEN_1566; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1568 = 8'h13 == _T_539 ? 8'h7d : _GEN_1567; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1569 = 8'h14 == _T_539 ? 8'hfa : _GEN_1568; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1570 = 8'h15 == _T_539 ? 8'h59 : _GEN_1569; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1571 = 8'h16 == _T_539 ? 8'h47 : _GEN_1570; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1572 = 8'h17 == _T_539 ? 8'hf0 : _GEN_1571; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1573 = 8'h18 == _T_539 ? 8'had : _GEN_1572; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1574 = 8'h19 == _T_539 ? 8'hd4 : _GEN_1573; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1575 = 8'h1a == _T_539 ? 8'ha2 : _GEN_1574; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1576 = 8'h1b == _T_539 ? 8'haf : _GEN_1575; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1577 = 8'h1c == _T_539 ? 8'h9c : _GEN_1576; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1578 = 8'h1d == _T_539 ? 8'ha4 : _GEN_1577; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1579 = 8'h1e == _T_539 ? 8'h72 : _GEN_1578; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1580 = 8'h1f == _T_539 ? 8'hc0 : _GEN_1579; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1581 = 8'h20 == _T_539 ? 8'hb7 : _GEN_1580; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1582 = 8'h21 == _T_539 ? 8'hfd : _GEN_1581; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1583 = 8'h22 == _T_539 ? 8'h93 : _GEN_1582; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1584 = 8'h23 == _T_539 ? 8'h26 : _GEN_1583; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1585 = 8'h24 == _T_539 ? 8'h36 : _GEN_1584; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1586 = 8'h25 == _T_539 ? 8'h3f : _GEN_1585; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1587 = 8'h26 == _T_539 ? 8'hf7 : _GEN_1586; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1588 = 8'h27 == _T_539 ? 8'hcc : _GEN_1587; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1589 = 8'h28 == _T_539 ? 8'h34 : _GEN_1588; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1590 = 8'h29 == _T_539 ? 8'ha5 : _GEN_1589; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1591 = 8'h2a == _T_539 ? 8'he5 : _GEN_1590; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1592 = 8'h2b == _T_539 ? 8'hf1 : _GEN_1591; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1593 = 8'h2c == _T_539 ? 8'h71 : _GEN_1592; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1594 = 8'h2d == _T_539 ? 8'hd8 : _GEN_1593; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1595 = 8'h2e == _T_539 ? 8'h31 : _GEN_1594; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1596 = 8'h2f == _T_539 ? 8'h15 : _GEN_1595; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1597 = 8'h30 == _T_539 ? 8'h4 : _GEN_1596; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1598 = 8'h31 == _T_539 ? 8'hc7 : _GEN_1597; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1599 = 8'h32 == _T_539 ? 8'h23 : _GEN_1598; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1600 = 8'h33 == _T_539 ? 8'hc3 : _GEN_1599; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1601 = 8'h34 == _T_539 ? 8'h18 : _GEN_1600; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1602 = 8'h35 == _T_539 ? 8'h96 : _GEN_1601; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1603 = 8'h36 == _T_539 ? 8'h5 : _GEN_1602; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1604 = 8'h37 == _T_539 ? 8'h9a : _GEN_1603; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1605 = 8'h38 == _T_539 ? 8'h7 : _GEN_1604; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1606 = 8'h39 == _T_539 ? 8'h12 : _GEN_1605; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1607 = 8'h3a == _T_539 ? 8'h80 : _GEN_1606; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1608 = 8'h3b == _T_539 ? 8'he2 : _GEN_1607; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1609 = 8'h3c == _T_539 ? 8'heb : _GEN_1608; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1610 = 8'h3d == _T_539 ? 8'h27 : _GEN_1609; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1611 = 8'h3e == _T_539 ? 8'hb2 : _GEN_1610; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1612 = 8'h3f == _T_539 ? 8'h75 : _GEN_1611; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1613 = 8'h40 == _T_539 ? 8'h9 : _GEN_1612; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1614 = 8'h41 == _T_539 ? 8'h83 : _GEN_1613; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1615 = 8'h42 == _T_539 ? 8'h2c : _GEN_1614; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1616 = 8'h43 == _T_539 ? 8'h1a : _GEN_1615; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1617 = 8'h44 == _T_539 ? 8'h1b : _GEN_1616; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1618 = 8'h45 == _T_539 ? 8'h6e : _GEN_1617; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1619 = 8'h46 == _T_539 ? 8'h5a : _GEN_1618; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1620 = 8'h47 == _T_539 ? 8'ha0 : _GEN_1619; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1621 = 8'h48 == _T_539 ? 8'h52 : _GEN_1620; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1622 = 8'h49 == _T_539 ? 8'h3b : _GEN_1621; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1623 = 8'h4a == _T_539 ? 8'hd6 : _GEN_1622; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1624 = 8'h4b == _T_539 ? 8'hb3 : _GEN_1623; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1625 = 8'h4c == _T_539 ? 8'h29 : _GEN_1624; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1626 = 8'h4d == _T_539 ? 8'he3 : _GEN_1625; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1627 = 8'h4e == _T_539 ? 8'h2f : _GEN_1626; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1628 = 8'h4f == _T_539 ? 8'h84 : _GEN_1627; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1629 = 8'h50 == _T_539 ? 8'h53 : _GEN_1628; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1630 = 8'h51 == _T_539 ? 8'hd1 : _GEN_1629; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1631 = 8'h52 == _T_539 ? 8'h0 : _GEN_1630; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1632 = 8'h53 == _T_539 ? 8'hed : _GEN_1631; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1633 = 8'h54 == _T_539 ? 8'h20 : _GEN_1632; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1634 = 8'h55 == _T_539 ? 8'hfc : _GEN_1633; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1635 = 8'h56 == _T_539 ? 8'hb1 : _GEN_1634; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1636 = 8'h57 == _T_539 ? 8'h5b : _GEN_1635; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1637 = 8'h58 == _T_539 ? 8'h6a : _GEN_1636; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1638 = 8'h59 == _T_539 ? 8'hcb : _GEN_1637; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1639 = 8'h5a == _T_539 ? 8'hbe : _GEN_1638; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1640 = 8'h5b == _T_539 ? 8'h39 : _GEN_1639; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1641 = 8'h5c == _T_539 ? 8'h4a : _GEN_1640; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1642 = 8'h5d == _T_539 ? 8'h4c : _GEN_1641; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1643 = 8'h5e == _T_539 ? 8'h58 : _GEN_1642; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1644 = 8'h5f == _T_539 ? 8'hcf : _GEN_1643; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1645 = 8'h60 == _T_539 ? 8'hd0 : _GEN_1644; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1646 = 8'h61 == _T_539 ? 8'hef : _GEN_1645; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1647 = 8'h62 == _T_539 ? 8'haa : _GEN_1646; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1648 = 8'h63 == _T_539 ? 8'hfb : _GEN_1647; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1649 = 8'h64 == _T_539 ? 8'h43 : _GEN_1648; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1650 = 8'h65 == _T_539 ? 8'h4d : _GEN_1649; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1651 = 8'h66 == _T_539 ? 8'h33 : _GEN_1650; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1652 = 8'h67 == _T_539 ? 8'h85 : _GEN_1651; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1653 = 8'h68 == _T_539 ? 8'h45 : _GEN_1652; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1654 = 8'h69 == _T_539 ? 8'hf9 : _GEN_1653; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1655 = 8'h6a == _T_539 ? 8'h2 : _GEN_1654; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1656 = 8'h6b == _T_539 ? 8'h7f : _GEN_1655; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1657 = 8'h6c == _T_539 ? 8'h50 : _GEN_1656; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1658 = 8'h6d == _T_539 ? 8'h3c : _GEN_1657; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1659 = 8'h6e == _T_539 ? 8'h9f : _GEN_1658; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1660 = 8'h6f == _T_539 ? 8'ha8 : _GEN_1659; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1661 = 8'h70 == _T_539 ? 8'h51 : _GEN_1660; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1662 = 8'h71 == _T_539 ? 8'ha3 : _GEN_1661; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1663 = 8'h72 == _T_539 ? 8'h40 : _GEN_1662; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1664 = 8'h73 == _T_539 ? 8'h8f : _GEN_1663; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1665 = 8'h74 == _T_539 ? 8'h92 : _GEN_1664; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1666 = 8'h75 == _T_539 ? 8'h9d : _GEN_1665; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1667 = 8'h76 == _T_539 ? 8'h38 : _GEN_1666; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1668 = 8'h77 == _T_539 ? 8'hf5 : _GEN_1667; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1669 = 8'h78 == _T_539 ? 8'hbc : _GEN_1668; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1670 = 8'h79 == _T_539 ? 8'hb6 : _GEN_1669; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1671 = 8'h7a == _T_539 ? 8'hda : _GEN_1670; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1672 = 8'h7b == _T_539 ? 8'h21 : _GEN_1671; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1673 = 8'h7c == _T_539 ? 8'h10 : _GEN_1672; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1674 = 8'h7d == _T_539 ? 8'hff : _GEN_1673; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1675 = 8'h7e == _T_539 ? 8'hf3 : _GEN_1674; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1676 = 8'h7f == _T_539 ? 8'hd2 : _GEN_1675; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1677 = 8'h80 == _T_539 ? 8'hcd : _GEN_1676; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1678 = 8'h81 == _T_539 ? 8'hc : _GEN_1677; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1679 = 8'h82 == _T_539 ? 8'h13 : _GEN_1678; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1680 = 8'h83 == _T_539 ? 8'hec : _GEN_1679; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1681 = 8'h84 == _T_539 ? 8'h5f : _GEN_1680; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1682 = 8'h85 == _T_539 ? 8'h97 : _GEN_1681; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1683 = 8'h86 == _T_539 ? 8'h44 : _GEN_1682; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1684 = 8'h87 == _T_539 ? 8'h17 : _GEN_1683; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1685 = 8'h88 == _T_539 ? 8'hc4 : _GEN_1684; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1686 = 8'h89 == _T_539 ? 8'ha7 : _GEN_1685; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1687 = 8'h8a == _T_539 ? 8'h7e : _GEN_1686; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1688 = 8'h8b == _T_539 ? 8'h3d : _GEN_1687; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1689 = 8'h8c == _T_539 ? 8'h64 : _GEN_1688; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1690 = 8'h8d == _T_539 ? 8'h5d : _GEN_1689; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1691 = 8'h8e == _T_539 ? 8'h19 : _GEN_1690; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1692 = 8'h8f == _T_539 ? 8'h73 : _GEN_1691; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1693 = 8'h90 == _T_539 ? 8'h60 : _GEN_1692; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1694 = 8'h91 == _T_539 ? 8'h81 : _GEN_1693; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1695 = 8'h92 == _T_539 ? 8'h4f : _GEN_1694; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1696 = 8'h93 == _T_539 ? 8'hdc : _GEN_1695; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1697 = 8'h94 == _T_539 ? 8'h22 : _GEN_1696; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1698 = 8'h95 == _T_539 ? 8'h2a : _GEN_1697; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1699 = 8'h96 == _T_539 ? 8'h90 : _GEN_1698; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1700 = 8'h97 == _T_539 ? 8'h88 : _GEN_1699; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1701 = 8'h98 == _T_539 ? 8'h46 : _GEN_1700; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1702 = 8'h99 == _T_539 ? 8'hee : _GEN_1701; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1703 = 8'h9a == _T_539 ? 8'hb8 : _GEN_1702; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1704 = 8'h9b == _T_539 ? 8'h14 : _GEN_1703; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1705 = 8'h9c == _T_539 ? 8'hde : _GEN_1704; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1706 = 8'h9d == _T_539 ? 8'h5e : _GEN_1705; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1707 = 8'h9e == _T_539 ? 8'hb : _GEN_1706; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1708 = 8'h9f == _T_539 ? 8'hdb : _GEN_1707; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1709 = 8'ha0 == _T_539 ? 8'he0 : _GEN_1708; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1710 = 8'ha1 == _T_539 ? 8'h32 : _GEN_1709; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1711 = 8'ha2 == _T_539 ? 8'h3a : _GEN_1710; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1712 = 8'ha3 == _T_539 ? 8'ha : _GEN_1711; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1713 = 8'ha4 == _T_539 ? 8'h49 : _GEN_1712; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1714 = 8'ha5 == _T_539 ? 8'h6 : _GEN_1713; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1715 = 8'ha6 == _T_539 ? 8'h24 : _GEN_1714; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1716 = 8'ha7 == _T_539 ? 8'h5c : _GEN_1715; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1717 = 8'ha8 == _T_539 ? 8'hc2 : _GEN_1716; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1718 = 8'ha9 == _T_539 ? 8'hd3 : _GEN_1717; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1719 = 8'haa == _T_539 ? 8'hac : _GEN_1718; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1720 = 8'hab == _T_539 ? 8'h62 : _GEN_1719; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1721 = 8'hac == _T_539 ? 8'h91 : _GEN_1720; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1722 = 8'had == _T_539 ? 8'h95 : _GEN_1721; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1723 = 8'hae == _T_539 ? 8'he4 : _GEN_1722; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1724 = 8'haf == _T_539 ? 8'h79 : _GEN_1723; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1725 = 8'hb0 == _T_539 ? 8'he7 : _GEN_1724; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1726 = 8'hb1 == _T_539 ? 8'hc8 : _GEN_1725; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1727 = 8'hb2 == _T_539 ? 8'h37 : _GEN_1726; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1728 = 8'hb3 == _T_539 ? 8'h6d : _GEN_1727; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1729 = 8'hb4 == _T_539 ? 8'h8d : _GEN_1728; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1730 = 8'hb5 == _T_539 ? 8'hd5 : _GEN_1729; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1731 = 8'hb6 == _T_539 ? 8'h4e : _GEN_1730; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1732 = 8'hb7 == _T_539 ? 8'ha9 : _GEN_1731; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1733 = 8'hb8 == _T_539 ? 8'h6c : _GEN_1732; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1734 = 8'hb9 == _T_539 ? 8'h56 : _GEN_1733; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1735 = 8'hba == _T_539 ? 8'hf4 : _GEN_1734; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1736 = 8'hbb == _T_539 ? 8'hea : _GEN_1735; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1737 = 8'hbc == _T_539 ? 8'h65 : _GEN_1736; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1738 = 8'hbd == _T_539 ? 8'h7a : _GEN_1737; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1739 = 8'hbe == _T_539 ? 8'hae : _GEN_1738; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1740 = 8'hbf == _T_539 ? 8'h8 : _GEN_1739; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1741 = 8'hc0 == _T_539 ? 8'hba : _GEN_1740; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1742 = 8'hc1 == _T_539 ? 8'h78 : _GEN_1741; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1743 = 8'hc2 == _T_539 ? 8'h25 : _GEN_1742; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1744 = 8'hc3 == _T_539 ? 8'h2e : _GEN_1743; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1745 = 8'hc4 == _T_539 ? 8'h1c : _GEN_1744; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1746 = 8'hc5 == _T_539 ? 8'ha6 : _GEN_1745; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1747 = 8'hc6 == _T_539 ? 8'hb4 : _GEN_1746; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1748 = 8'hc7 == _T_539 ? 8'hc6 : _GEN_1747; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1749 = 8'hc8 == _T_539 ? 8'he8 : _GEN_1748; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1750 = 8'hc9 == _T_539 ? 8'hdd : _GEN_1749; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1751 = 8'hca == _T_539 ? 8'h74 : _GEN_1750; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1752 = 8'hcb == _T_539 ? 8'h1f : _GEN_1751; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1753 = 8'hcc == _T_539 ? 8'h4b : _GEN_1752; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1754 = 8'hcd == _T_539 ? 8'hbd : _GEN_1753; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1755 = 8'hce == _T_539 ? 8'h8b : _GEN_1754; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1756 = 8'hcf == _T_539 ? 8'h8a : _GEN_1755; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1757 = 8'hd0 == _T_539 ? 8'h70 : _GEN_1756; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1758 = 8'hd1 == _T_539 ? 8'h3e : _GEN_1757; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1759 = 8'hd2 == _T_539 ? 8'hb5 : _GEN_1758; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1760 = 8'hd3 == _T_539 ? 8'h66 : _GEN_1759; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1761 = 8'hd4 == _T_539 ? 8'h48 : _GEN_1760; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1762 = 8'hd5 == _T_539 ? 8'h3 : _GEN_1761; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1763 = 8'hd6 == _T_539 ? 8'hf6 : _GEN_1762; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1764 = 8'hd7 == _T_539 ? 8'he : _GEN_1763; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1765 = 8'hd8 == _T_539 ? 8'h61 : _GEN_1764; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1766 = 8'hd9 == _T_539 ? 8'h35 : _GEN_1765; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1767 = 8'hda == _T_539 ? 8'h57 : _GEN_1766; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1768 = 8'hdb == _T_539 ? 8'hb9 : _GEN_1767; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1769 = 8'hdc == _T_539 ? 8'h86 : _GEN_1768; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1770 = 8'hdd == _T_539 ? 8'hc1 : _GEN_1769; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1771 = 8'hde == _T_539 ? 8'h1d : _GEN_1770; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1772 = 8'hdf == _T_539 ? 8'h9e : _GEN_1771; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1773 = 8'he0 == _T_539 ? 8'he1 : _GEN_1772; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1774 = 8'he1 == _T_539 ? 8'hf8 : _GEN_1773; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1775 = 8'he2 == _T_539 ? 8'h98 : _GEN_1774; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1776 = 8'he3 == _T_539 ? 8'h11 : _GEN_1775; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1777 = 8'he4 == _T_539 ? 8'h69 : _GEN_1776; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1778 = 8'he5 == _T_539 ? 8'hd9 : _GEN_1777; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1779 = 8'he6 == _T_539 ? 8'h8e : _GEN_1778; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1780 = 8'he7 == _T_539 ? 8'h94 : _GEN_1779; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1781 = 8'he8 == _T_539 ? 8'h9b : _GEN_1780; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1782 = 8'he9 == _T_539 ? 8'h1e : _GEN_1781; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1783 = 8'hea == _T_539 ? 8'h87 : _GEN_1782; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1784 = 8'heb == _T_539 ? 8'he9 : _GEN_1783; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1785 = 8'hec == _T_539 ? 8'hce : _GEN_1784; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1786 = 8'hed == _T_539 ? 8'h55 : _GEN_1785; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1787 = 8'hee == _T_539 ? 8'h28 : _GEN_1786; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1788 = 8'hef == _T_539 ? 8'hdf : _GEN_1787; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1789 = 8'hf0 == _T_539 ? 8'h8c : _GEN_1788; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1790 = 8'hf1 == _T_539 ? 8'ha1 : _GEN_1789; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1791 = 8'hf2 == _T_539 ? 8'h89 : _GEN_1790; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1792 = 8'hf3 == _T_539 ? 8'hd : _GEN_1791; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1793 = 8'hf4 == _T_539 ? 8'hbf : _GEN_1792; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1794 = 8'hf5 == _T_539 ? 8'he6 : _GEN_1793; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1795 = 8'hf6 == _T_539 ? 8'h42 : _GEN_1794; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1796 = 8'hf7 == _T_539 ? 8'h68 : _GEN_1795; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1797 = 8'hf8 == _T_539 ? 8'h41 : _GEN_1796; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1798 = 8'hf9 == _T_539 ? 8'h99 : _GEN_1797; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1799 = 8'hfa == _T_539 ? 8'h2d : _GEN_1798; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1800 = 8'hfb == _T_539 ? 8'hf : _GEN_1799; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1801 = 8'hfc == _T_539 ? 8'hb0 : _GEN_1800; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1802 = 8'hfd == _T_539 ? 8'h54 : _GEN_1801; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1803 = 8'hfe == _T_539 ? 8'hbb : _GEN_1802; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1804 = 8'hff == _T_539 ? 8'h16 : _GEN_1803; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1805 = 8'h1 == _T_537 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1806 = 8'h2 == _T_537 ? 8'h77 : _GEN_1805; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1807 = 8'h3 == _T_537 ? 8'h7b : _GEN_1806; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1808 = 8'h4 == _T_537 ? 8'hf2 : _GEN_1807; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1809 = 8'h5 == _T_537 ? 8'h6b : _GEN_1808; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1810 = 8'h6 == _T_537 ? 8'h6f : _GEN_1809; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1811 = 8'h7 == _T_537 ? 8'hc5 : _GEN_1810; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1812 = 8'h8 == _T_537 ? 8'h30 : _GEN_1811; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1813 = 8'h9 == _T_537 ? 8'h1 : _GEN_1812; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1814 = 8'ha == _T_537 ? 8'h67 : _GEN_1813; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1815 = 8'hb == _T_537 ? 8'h2b : _GEN_1814; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1816 = 8'hc == _T_537 ? 8'hfe : _GEN_1815; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1817 = 8'hd == _T_537 ? 8'hd7 : _GEN_1816; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1818 = 8'he == _T_537 ? 8'hab : _GEN_1817; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1819 = 8'hf == _T_537 ? 8'h76 : _GEN_1818; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1820 = 8'h10 == _T_537 ? 8'hca : _GEN_1819; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1821 = 8'h11 == _T_537 ? 8'h82 : _GEN_1820; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1822 = 8'h12 == _T_537 ? 8'hc9 : _GEN_1821; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1823 = 8'h13 == _T_537 ? 8'h7d : _GEN_1822; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1824 = 8'h14 == _T_537 ? 8'hfa : _GEN_1823; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1825 = 8'h15 == _T_537 ? 8'h59 : _GEN_1824; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1826 = 8'h16 == _T_537 ? 8'h47 : _GEN_1825; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1827 = 8'h17 == _T_537 ? 8'hf0 : _GEN_1826; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1828 = 8'h18 == _T_537 ? 8'had : _GEN_1827; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1829 = 8'h19 == _T_537 ? 8'hd4 : _GEN_1828; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1830 = 8'h1a == _T_537 ? 8'ha2 : _GEN_1829; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1831 = 8'h1b == _T_537 ? 8'haf : _GEN_1830; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1832 = 8'h1c == _T_537 ? 8'h9c : _GEN_1831; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1833 = 8'h1d == _T_537 ? 8'ha4 : _GEN_1832; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1834 = 8'h1e == _T_537 ? 8'h72 : _GEN_1833; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1835 = 8'h1f == _T_537 ? 8'hc0 : _GEN_1834; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1836 = 8'h20 == _T_537 ? 8'hb7 : _GEN_1835; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1837 = 8'h21 == _T_537 ? 8'hfd : _GEN_1836; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1838 = 8'h22 == _T_537 ? 8'h93 : _GEN_1837; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1839 = 8'h23 == _T_537 ? 8'h26 : _GEN_1838; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1840 = 8'h24 == _T_537 ? 8'h36 : _GEN_1839; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1841 = 8'h25 == _T_537 ? 8'h3f : _GEN_1840; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1842 = 8'h26 == _T_537 ? 8'hf7 : _GEN_1841; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1843 = 8'h27 == _T_537 ? 8'hcc : _GEN_1842; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1844 = 8'h28 == _T_537 ? 8'h34 : _GEN_1843; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1845 = 8'h29 == _T_537 ? 8'ha5 : _GEN_1844; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1846 = 8'h2a == _T_537 ? 8'he5 : _GEN_1845; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1847 = 8'h2b == _T_537 ? 8'hf1 : _GEN_1846; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1848 = 8'h2c == _T_537 ? 8'h71 : _GEN_1847; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1849 = 8'h2d == _T_537 ? 8'hd8 : _GEN_1848; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1850 = 8'h2e == _T_537 ? 8'h31 : _GEN_1849; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1851 = 8'h2f == _T_537 ? 8'h15 : _GEN_1850; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1852 = 8'h30 == _T_537 ? 8'h4 : _GEN_1851; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1853 = 8'h31 == _T_537 ? 8'hc7 : _GEN_1852; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1854 = 8'h32 == _T_537 ? 8'h23 : _GEN_1853; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1855 = 8'h33 == _T_537 ? 8'hc3 : _GEN_1854; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1856 = 8'h34 == _T_537 ? 8'h18 : _GEN_1855; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1857 = 8'h35 == _T_537 ? 8'h96 : _GEN_1856; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1858 = 8'h36 == _T_537 ? 8'h5 : _GEN_1857; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1859 = 8'h37 == _T_537 ? 8'h9a : _GEN_1858; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1860 = 8'h38 == _T_537 ? 8'h7 : _GEN_1859; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1861 = 8'h39 == _T_537 ? 8'h12 : _GEN_1860; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1862 = 8'h3a == _T_537 ? 8'h80 : _GEN_1861; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1863 = 8'h3b == _T_537 ? 8'he2 : _GEN_1862; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1864 = 8'h3c == _T_537 ? 8'heb : _GEN_1863; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1865 = 8'h3d == _T_537 ? 8'h27 : _GEN_1864; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1866 = 8'h3e == _T_537 ? 8'hb2 : _GEN_1865; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1867 = 8'h3f == _T_537 ? 8'h75 : _GEN_1866; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1868 = 8'h40 == _T_537 ? 8'h9 : _GEN_1867; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1869 = 8'h41 == _T_537 ? 8'h83 : _GEN_1868; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1870 = 8'h42 == _T_537 ? 8'h2c : _GEN_1869; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1871 = 8'h43 == _T_537 ? 8'h1a : _GEN_1870; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1872 = 8'h44 == _T_537 ? 8'h1b : _GEN_1871; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1873 = 8'h45 == _T_537 ? 8'h6e : _GEN_1872; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1874 = 8'h46 == _T_537 ? 8'h5a : _GEN_1873; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1875 = 8'h47 == _T_537 ? 8'ha0 : _GEN_1874; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1876 = 8'h48 == _T_537 ? 8'h52 : _GEN_1875; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1877 = 8'h49 == _T_537 ? 8'h3b : _GEN_1876; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1878 = 8'h4a == _T_537 ? 8'hd6 : _GEN_1877; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1879 = 8'h4b == _T_537 ? 8'hb3 : _GEN_1878; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1880 = 8'h4c == _T_537 ? 8'h29 : _GEN_1879; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1881 = 8'h4d == _T_537 ? 8'he3 : _GEN_1880; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1882 = 8'h4e == _T_537 ? 8'h2f : _GEN_1881; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1883 = 8'h4f == _T_537 ? 8'h84 : _GEN_1882; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1884 = 8'h50 == _T_537 ? 8'h53 : _GEN_1883; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1885 = 8'h51 == _T_537 ? 8'hd1 : _GEN_1884; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1886 = 8'h52 == _T_537 ? 8'h0 : _GEN_1885; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1887 = 8'h53 == _T_537 ? 8'hed : _GEN_1886; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1888 = 8'h54 == _T_537 ? 8'h20 : _GEN_1887; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1889 = 8'h55 == _T_537 ? 8'hfc : _GEN_1888; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1890 = 8'h56 == _T_537 ? 8'hb1 : _GEN_1889; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1891 = 8'h57 == _T_537 ? 8'h5b : _GEN_1890; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1892 = 8'h58 == _T_537 ? 8'h6a : _GEN_1891; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1893 = 8'h59 == _T_537 ? 8'hcb : _GEN_1892; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1894 = 8'h5a == _T_537 ? 8'hbe : _GEN_1893; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1895 = 8'h5b == _T_537 ? 8'h39 : _GEN_1894; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1896 = 8'h5c == _T_537 ? 8'h4a : _GEN_1895; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1897 = 8'h5d == _T_537 ? 8'h4c : _GEN_1896; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1898 = 8'h5e == _T_537 ? 8'h58 : _GEN_1897; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1899 = 8'h5f == _T_537 ? 8'hcf : _GEN_1898; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1900 = 8'h60 == _T_537 ? 8'hd0 : _GEN_1899; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1901 = 8'h61 == _T_537 ? 8'hef : _GEN_1900; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1902 = 8'h62 == _T_537 ? 8'haa : _GEN_1901; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1903 = 8'h63 == _T_537 ? 8'hfb : _GEN_1902; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1904 = 8'h64 == _T_537 ? 8'h43 : _GEN_1903; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1905 = 8'h65 == _T_537 ? 8'h4d : _GEN_1904; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1906 = 8'h66 == _T_537 ? 8'h33 : _GEN_1905; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1907 = 8'h67 == _T_537 ? 8'h85 : _GEN_1906; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1908 = 8'h68 == _T_537 ? 8'h45 : _GEN_1907; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1909 = 8'h69 == _T_537 ? 8'hf9 : _GEN_1908; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1910 = 8'h6a == _T_537 ? 8'h2 : _GEN_1909; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1911 = 8'h6b == _T_537 ? 8'h7f : _GEN_1910; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1912 = 8'h6c == _T_537 ? 8'h50 : _GEN_1911; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1913 = 8'h6d == _T_537 ? 8'h3c : _GEN_1912; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1914 = 8'h6e == _T_537 ? 8'h9f : _GEN_1913; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1915 = 8'h6f == _T_537 ? 8'ha8 : _GEN_1914; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1916 = 8'h70 == _T_537 ? 8'h51 : _GEN_1915; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1917 = 8'h71 == _T_537 ? 8'ha3 : _GEN_1916; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1918 = 8'h72 == _T_537 ? 8'h40 : _GEN_1917; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1919 = 8'h73 == _T_537 ? 8'h8f : _GEN_1918; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1920 = 8'h74 == _T_537 ? 8'h92 : _GEN_1919; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1921 = 8'h75 == _T_537 ? 8'h9d : _GEN_1920; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1922 = 8'h76 == _T_537 ? 8'h38 : _GEN_1921; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1923 = 8'h77 == _T_537 ? 8'hf5 : _GEN_1922; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1924 = 8'h78 == _T_537 ? 8'hbc : _GEN_1923; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1925 = 8'h79 == _T_537 ? 8'hb6 : _GEN_1924; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1926 = 8'h7a == _T_537 ? 8'hda : _GEN_1925; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1927 = 8'h7b == _T_537 ? 8'h21 : _GEN_1926; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1928 = 8'h7c == _T_537 ? 8'h10 : _GEN_1927; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1929 = 8'h7d == _T_537 ? 8'hff : _GEN_1928; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1930 = 8'h7e == _T_537 ? 8'hf3 : _GEN_1929; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1931 = 8'h7f == _T_537 ? 8'hd2 : _GEN_1930; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1932 = 8'h80 == _T_537 ? 8'hcd : _GEN_1931; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1933 = 8'h81 == _T_537 ? 8'hc : _GEN_1932; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1934 = 8'h82 == _T_537 ? 8'h13 : _GEN_1933; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1935 = 8'h83 == _T_537 ? 8'hec : _GEN_1934; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1936 = 8'h84 == _T_537 ? 8'h5f : _GEN_1935; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1937 = 8'h85 == _T_537 ? 8'h97 : _GEN_1936; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1938 = 8'h86 == _T_537 ? 8'h44 : _GEN_1937; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1939 = 8'h87 == _T_537 ? 8'h17 : _GEN_1938; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1940 = 8'h88 == _T_537 ? 8'hc4 : _GEN_1939; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1941 = 8'h89 == _T_537 ? 8'ha7 : _GEN_1940; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1942 = 8'h8a == _T_537 ? 8'h7e : _GEN_1941; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1943 = 8'h8b == _T_537 ? 8'h3d : _GEN_1942; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1944 = 8'h8c == _T_537 ? 8'h64 : _GEN_1943; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1945 = 8'h8d == _T_537 ? 8'h5d : _GEN_1944; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1946 = 8'h8e == _T_537 ? 8'h19 : _GEN_1945; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1947 = 8'h8f == _T_537 ? 8'h73 : _GEN_1946; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1948 = 8'h90 == _T_537 ? 8'h60 : _GEN_1947; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1949 = 8'h91 == _T_537 ? 8'h81 : _GEN_1948; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1950 = 8'h92 == _T_537 ? 8'h4f : _GEN_1949; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1951 = 8'h93 == _T_537 ? 8'hdc : _GEN_1950; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1952 = 8'h94 == _T_537 ? 8'h22 : _GEN_1951; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1953 = 8'h95 == _T_537 ? 8'h2a : _GEN_1952; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1954 = 8'h96 == _T_537 ? 8'h90 : _GEN_1953; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1955 = 8'h97 == _T_537 ? 8'h88 : _GEN_1954; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1956 = 8'h98 == _T_537 ? 8'h46 : _GEN_1955; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1957 = 8'h99 == _T_537 ? 8'hee : _GEN_1956; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1958 = 8'h9a == _T_537 ? 8'hb8 : _GEN_1957; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1959 = 8'h9b == _T_537 ? 8'h14 : _GEN_1958; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1960 = 8'h9c == _T_537 ? 8'hde : _GEN_1959; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1961 = 8'h9d == _T_537 ? 8'h5e : _GEN_1960; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1962 = 8'h9e == _T_537 ? 8'hb : _GEN_1961; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1963 = 8'h9f == _T_537 ? 8'hdb : _GEN_1962; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1964 = 8'ha0 == _T_537 ? 8'he0 : _GEN_1963; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1965 = 8'ha1 == _T_537 ? 8'h32 : _GEN_1964; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1966 = 8'ha2 == _T_537 ? 8'h3a : _GEN_1965; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1967 = 8'ha3 == _T_537 ? 8'ha : _GEN_1966; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1968 = 8'ha4 == _T_537 ? 8'h49 : _GEN_1967; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1969 = 8'ha5 == _T_537 ? 8'h6 : _GEN_1968; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1970 = 8'ha6 == _T_537 ? 8'h24 : _GEN_1969; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1971 = 8'ha7 == _T_537 ? 8'h5c : _GEN_1970; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1972 = 8'ha8 == _T_537 ? 8'hc2 : _GEN_1971; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1973 = 8'ha9 == _T_537 ? 8'hd3 : _GEN_1972; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1974 = 8'haa == _T_537 ? 8'hac : _GEN_1973; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1975 = 8'hab == _T_537 ? 8'h62 : _GEN_1974; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1976 = 8'hac == _T_537 ? 8'h91 : _GEN_1975; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1977 = 8'had == _T_537 ? 8'h95 : _GEN_1976; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1978 = 8'hae == _T_537 ? 8'he4 : _GEN_1977; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1979 = 8'haf == _T_537 ? 8'h79 : _GEN_1978; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1980 = 8'hb0 == _T_537 ? 8'he7 : _GEN_1979; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1981 = 8'hb1 == _T_537 ? 8'hc8 : _GEN_1980; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1982 = 8'hb2 == _T_537 ? 8'h37 : _GEN_1981; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1983 = 8'hb3 == _T_537 ? 8'h6d : _GEN_1982; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1984 = 8'hb4 == _T_537 ? 8'h8d : _GEN_1983; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1985 = 8'hb5 == _T_537 ? 8'hd5 : _GEN_1984; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1986 = 8'hb6 == _T_537 ? 8'h4e : _GEN_1985; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1987 = 8'hb7 == _T_537 ? 8'ha9 : _GEN_1986; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1988 = 8'hb8 == _T_537 ? 8'h6c : _GEN_1987; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1989 = 8'hb9 == _T_537 ? 8'h56 : _GEN_1988; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1990 = 8'hba == _T_537 ? 8'hf4 : _GEN_1989; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1991 = 8'hbb == _T_537 ? 8'hea : _GEN_1990; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1992 = 8'hbc == _T_537 ? 8'h65 : _GEN_1991; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1993 = 8'hbd == _T_537 ? 8'h7a : _GEN_1992; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1994 = 8'hbe == _T_537 ? 8'hae : _GEN_1993; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1995 = 8'hbf == _T_537 ? 8'h8 : _GEN_1994; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1996 = 8'hc0 == _T_537 ? 8'hba : _GEN_1995; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1997 = 8'hc1 == _T_537 ? 8'h78 : _GEN_1996; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1998 = 8'hc2 == _T_537 ? 8'h25 : _GEN_1997; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_1999 = 8'hc3 == _T_537 ? 8'h2e : _GEN_1998; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2000 = 8'hc4 == _T_537 ? 8'h1c : _GEN_1999; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2001 = 8'hc5 == _T_537 ? 8'ha6 : _GEN_2000; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2002 = 8'hc6 == _T_537 ? 8'hb4 : _GEN_2001; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2003 = 8'hc7 == _T_537 ? 8'hc6 : _GEN_2002; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2004 = 8'hc8 == _T_537 ? 8'he8 : _GEN_2003; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2005 = 8'hc9 == _T_537 ? 8'hdd : _GEN_2004; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2006 = 8'hca == _T_537 ? 8'h74 : _GEN_2005; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2007 = 8'hcb == _T_537 ? 8'h1f : _GEN_2006; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2008 = 8'hcc == _T_537 ? 8'h4b : _GEN_2007; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2009 = 8'hcd == _T_537 ? 8'hbd : _GEN_2008; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2010 = 8'hce == _T_537 ? 8'h8b : _GEN_2009; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2011 = 8'hcf == _T_537 ? 8'h8a : _GEN_2010; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2012 = 8'hd0 == _T_537 ? 8'h70 : _GEN_2011; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2013 = 8'hd1 == _T_537 ? 8'h3e : _GEN_2012; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2014 = 8'hd2 == _T_537 ? 8'hb5 : _GEN_2013; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2015 = 8'hd3 == _T_537 ? 8'h66 : _GEN_2014; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2016 = 8'hd4 == _T_537 ? 8'h48 : _GEN_2015; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2017 = 8'hd5 == _T_537 ? 8'h3 : _GEN_2016; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2018 = 8'hd6 == _T_537 ? 8'hf6 : _GEN_2017; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2019 = 8'hd7 == _T_537 ? 8'he : _GEN_2018; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2020 = 8'hd8 == _T_537 ? 8'h61 : _GEN_2019; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2021 = 8'hd9 == _T_537 ? 8'h35 : _GEN_2020; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2022 = 8'hda == _T_537 ? 8'h57 : _GEN_2021; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2023 = 8'hdb == _T_537 ? 8'hb9 : _GEN_2022; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2024 = 8'hdc == _T_537 ? 8'h86 : _GEN_2023; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2025 = 8'hdd == _T_537 ? 8'hc1 : _GEN_2024; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2026 = 8'hde == _T_537 ? 8'h1d : _GEN_2025; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2027 = 8'hdf == _T_537 ? 8'h9e : _GEN_2026; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2028 = 8'he0 == _T_537 ? 8'he1 : _GEN_2027; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2029 = 8'he1 == _T_537 ? 8'hf8 : _GEN_2028; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2030 = 8'he2 == _T_537 ? 8'h98 : _GEN_2029; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2031 = 8'he3 == _T_537 ? 8'h11 : _GEN_2030; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2032 = 8'he4 == _T_537 ? 8'h69 : _GEN_2031; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2033 = 8'he5 == _T_537 ? 8'hd9 : _GEN_2032; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2034 = 8'he6 == _T_537 ? 8'h8e : _GEN_2033; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2035 = 8'he7 == _T_537 ? 8'h94 : _GEN_2034; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2036 = 8'he8 == _T_537 ? 8'h9b : _GEN_2035; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2037 = 8'he9 == _T_537 ? 8'h1e : _GEN_2036; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2038 = 8'hea == _T_537 ? 8'h87 : _GEN_2037; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2039 = 8'heb == _T_537 ? 8'he9 : _GEN_2038; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2040 = 8'hec == _T_537 ? 8'hce : _GEN_2039; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2041 = 8'hed == _T_537 ? 8'h55 : _GEN_2040; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2042 = 8'hee == _T_537 ? 8'h28 : _GEN_2041; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2043 = 8'hef == _T_537 ? 8'hdf : _GEN_2042; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2044 = 8'hf0 == _T_537 ? 8'h8c : _GEN_2043; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2045 = 8'hf1 == _T_537 ? 8'ha1 : _GEN_2044; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2046 = 8'hf2 == _T_537 ? 8'h89 : _GEN_2045; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2047 = 8'hf3 == _T_537 ? 8'hd : _GEN_2046; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2048 = 8'hf4 == _T_537 ? 8'hbf : _GEN_2047; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2049 = 8'hf5 == _T_537 ? 8'he6 : _GEN_2048; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2050 = 8'hf6 == _T_537 ? 8'h42 : _GEN_2049; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2051 = 8'hf7 == _T_537 ? 8'h68 : _GEN_2050; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2052 = 8'hf8 == _T_537 ? 8'h41 : _GEN_2051; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2053 = 8'hf9 == _T_537 ? 8'h99 : _GEN_2052; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2054 = 8'hfa == _T_537 ? 8'h2d : _GEN_2053; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2055 = 8'hfb == _T_537 ? 8'hf : _GEN_2054; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2056 = 8'hfc == _T_537 ? 8'hb0 : _GEN_2055; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2057 = 8'hfd == _T_537 ? 8'h54 : _GEN_2056; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2058 = 8'hfe == _T_537 ? 8'hbb : _GEN_2057; // @[Cat.scala 30:58:@2074.4]
  assign _GEN_2059 = 8'hff == _T_537 ? 8'h16 : _GEN_2058; // @[Cat.scala 30:58:@2074.4]
  assign _T_542 = {_GEN_1804,_GEN_2059}; // @[Cat.scala 30:58:@2074.4]
  assign x1 = {_T_542,_T_541}; // @[Cat.scala 30:58:@2075.4]
  assign _T_543 = io_addr2[39:32]; // @[sbox.scala 62:25:@2076.4]
  assign _T_545 = io_addr2[47:40]; // @[sbox.scala 63:25:@2077.4]
  assign _T_547 = io_addr2[55:48]; // @[sbox.scala 64:26:@2078.4]
  assign _T_549 = io_addr2[63:56]; // @[sbox.scala 65:26:@2079.4]
  assign _GEN_2060 = 8'h1 == _T_545 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2061 = 8'h2 == _T_545 ? 8'h77 : _GEN_2060; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2062 = 8'h3 == _T_545 ? 8'h7b : _GEN_2061; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2063 = 8'h4 == _T_545 ? 8'hf2 : _GEN_2062; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2064 = 8'h5 == _T_545 ? 8'h6b : _GEN_2063; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2065 = 8'h6 == _T_545 ? 8'h6f : _GEN_2064; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2066 = 8'h7 == _T_545 ? 8'hc5 : _GEN_2065; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2067 = 8'h8 == _T_545 ? 8'h30 : _GEN_2066; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2068 = 8'h9 == _T_545 ? 8'h1 : _GEN_2067; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2069 = 8'ha == _T_545 ? 8'h67 : _GEN_2068; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2070 = 8'hb == _T_545 ? 8'h2b : _GEN_2069; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2071 = 8'hc == _T_545 ? 8'hfe : _GEN_2070; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2072 = 8'hd == _T_545 ? 8'hd7 : _GEN_2071; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2073 = 8'he == _T_545 ? 8'hab : _GEN_2072; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2074 = 8'hf == _T_545 ? 8'h76 : _GEN_2073; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2075 = 8'h10 == _T_545 ? 8'hca : _GEN_2074; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2076 = 8'h11 == _T_545 ? 8'h82 : _GEN_2075; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2077 = 8'h12 == _T_545 ? 8'hc9 : _GEN_2076; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2078 = 8'h13 == _T_545 ? 8'h7d : _GEN_2077; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2079 = 8'h14 == _T_545 ? 8'hfa : _GEN_2078; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2080 = 8'h15 == _T_545 ? 8'h59 : _GEN_2079; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2081 = 8'h16 == _T_545 ? 8'h47 : _GEN_2080; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2082 = 8'h17 == _T_545 ? 8'hf0 : _GEN_2081; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2083 = 8'h18 == _T_545 ? 8'had : _GEN_2082; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2084 = 8'h19 == _T_545 ? 8'hd4 : _GEN_2083; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2085 = 8'h1a == _T_545 ? 8'ha2 : _GEN_2084; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2086 = 8'h1b == _T_545 ? 8'haf : _GEN_2085; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2087 = 8'h1c == _T_545 ? 8'h9c : _GEN_2086; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2088 = 8'h1d == _T_545 ? 8'ha4 : _GEN_2087; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2089 = 8'h1e == _T_545 ? 8'h72 : _GEN_2088; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2090 = 8'h1f == _T_545 ? 8'hc0 : _GEN_2089; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2091 = 8'h20 == _T_545 ? 8'hb7 : _GEN_2090; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2092 = 8'h21 == _T_545 ? 8'hfd : _GEN_2091; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2093 = 8'h22 == _T_545 ? 8'h93 : _GEN_2092; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2094 = 8'h23 == _T_545 ? 8'h26 : _GEN_2093; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2095 = 8'h24 == _T_545 ? 8'h36 : _GEN_2094; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2096 = 8'h25 == _T_545 ? 8'h3f : _GEN_2095; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2097 = 8'h26 == _T_545 ? 8'hf7 : _GEN_2096; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2098 = 8'h27 == _T_545 ? 8'hcc : _GEN_2097; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2099 = 8'h28 == _T_545 ? 8'h34 : _GEN_2098; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2100 = 8'h29 == _T_545 ? 8'ha5 : _GEN_2099; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2101 = 8'h2a == _T_545 ? 8'he5 : _GEN_2100; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2102 = 8'h2b == _T_545 ? 8'hf1 : _GEN_2101; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2103 = 8'h2c == _T_545 ? 8'h71 : _GEN_2102; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2104 = 8'h2d == _T_545 ? 8'hd8 : _GEN_2103; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2105 = 8'h2e == _T_545 ? 8'h31 : _GEN_2104; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2106 = 8'h2f == _T_545 ? 8'h15 : _GEN_2105; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2107 = 8'h30 == _T_545 ? 8'h4 : _GEN_2106; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2108 = 8'h31 == _T_545 ? 8'hc7 : _GEN_2107; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2109 = 8'h32 == _T_545 ? 8'h23 : _GEN_2108; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2110 = 8'h33 == _T_545 ? 8'hc3 : _GEN_2109; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2111 = 8'h34 == _T_545 ? 8'h18 : _GEN_2110; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2112 = 8'h35 == _T_545 ? 8'h96 : _GEN_2111; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2113 = 8'h36 == _T_545 ? 8'h5 : _GEN_2112; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2114 = 8'h37 == _T_545 ? 8'h9a : _GEN_2113; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2115 = 8'h38 == _T_545 ? 8'h7 : _GEN_2114; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2116 = 8'h39 == _T_545 ? 8'h12 : _GEN_2115; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2117 = 8'h3a == _T_545 ? 8'h80 : _GEN_2116; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2118 = 8'h3b == _T_545 ? 8'he2 : _GEN_2117; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2119 = 8'h3c == _T_545 ? 8'heb : _GEN_2118; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2120 = 8'h3d == _T_545 ? 8'h27 : _GEN_2119; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2121 = 8'h3e == _T_545 ? 8'hb2 : _GEN_2120; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2122 = 8'h3f == _T_545 ? 8'h75 : _GEN_2121; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2123 = 8'h40 == _T_545 ? 8'h9 : _GEN_2122; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2124 = 8'h41 == _T_545 ? 8'h83 : _GEN_2123; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2125 = 8'h42 == _T_545 ? 8'h2c : _GEN_2124; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2126 = 8'h43 == _T_545 ? 8'h1a : _GEN_2125; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2127 = 8'h44 == _T_545 ? 8'h1b : _GEN_2126; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2128 = 8'h45 == _T_545 ? 8'h6e : _GEN_2127; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2129 = 8'h46 == _T_545 ? 8'h5a : _GEN_2128; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2130 = 8'h47 == _T_545 ? 8'ha0 : _GEN_2129; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2131 = 8'h48 == _T_545 ? 8'h52 : _GEN_2130; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2132 = 8'h49 == _T_545 ? 8'h3b : _GEN_2131; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2133 = 8'h4a == _T_545 ? 8'hd6 : _GEN_2132; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2134 = 8'h4b == _T_545 ? 8'hb3 : _GEN_2133; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2135 = 8'h4c == _T_545 ? 8'h29 : _GEN_2134; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2136 = 8'h4d == _T_545 ? 8'he3 : _GEN_2135; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2137 = 8'h4e == _T_545 ? 8'h2f : _GEN_2136; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2138 = 8'h4f == _T_545 ? 8'h84 : _GEN_2137; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2139 = 8'h50 == _T_545 ? 8'h53 : _GEN_2138; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2140 = 8'h51 == _T_545 ? 8'hd1 : _GEN_2139; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2141 = 8'h52 == _T_545 ? 8'h0 : _GEN_2140; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2142 = 8'h53 == _T_545 ? 8'hed : _GEN_2141; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2143 = 8'h54 == _T_545 ? 8'h20 : _GEN_2142; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2144 = 8'h55 == _T_545 ? 8'hfc : _GEN_2143; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2145 = 8'h56 == _T_545 ? 8'hb1 : _GEN_2144; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2146 = 8'h57 == _T_545 ? 8'h5b : _GEN_2145; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2147 = 8'h58 == _T_545 ? 8'h6a : _GEN_2146; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2148 = 8'h59 == _T_545 ? 8'hcb : _GEN_2147; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2149 = 8'h5a == _T_545 ? 8'hbe : _GEN_2148; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2150 = 8'h5b == _T_545 ? 8'h39 : _GEN_2149; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2151 = 8'h5c == _T_545 ? 8'h4a : _GEN_2150; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2152 = 8'h5d == _T_545 ? 8'h4c : _GEN_2151; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2153 = 8'h5e == _T_545 ? 8'h58 : _GEN_2152; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2154 = 8'h5f == _T_545 ? 8'hcf : _GEN_2153; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2155 = 8'h60 == _T_545 ? 8'hd0 : _GEN_2154; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2156 = 8'h61 == _T_545 ? 8'hef : _GEN_2155; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2157 = 8'h62 == _T_545 ? 8'haa : _GEN_2156; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2158 = 8'h63 == _T_545 ? 8'hfb : _GEN_2157; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2159 = 8'h64 == _T_545 ? 8'h43 : _GEN_2158; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2160 = 8'h65 == _T_545 ? 8'h4d : _GEN_2159; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2161 = 8'h66 == _T_545 ? 8'h33 : _GEN_2160; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2162 = 8'h67 == _T_545 ? 8'h85 : _GEN_2161; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2163 = 8'h68 == _T_545 ? 8'h45 : _GEN_2162; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2164 = 8'h69 == _T_545 ? 8'hf9 : _GEN_2163; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2165 = 8'h6a == _T_545 ? 8'h2 : _GEN_2164; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2166 = 8'h6b == _T_545 ? 8'h7f : _GEN_2165; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2167 = 8'h6c == _T_545 ? 8'h50 : _GEN_2166; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2168 = 8'h6d == _T_545 ? 8'h3c : _GEN_2167; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2169 = 8'h6e == _T_545 ? 8'h9f : _GEN_2168; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2170 = 8'h6f == _T_545 ? 8'ha8 : _GEN_2169; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2171 = 8'h70 == _T_545 ? 8'h51 : _GEN_2170; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2172 = 8'h71 == _T_545 ? 8'ha3 : _GEN_2171; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2173 = 8'h72 == _T_545 ? 8'h40 : _GEN_2172; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2174 = 8'h73 == _T_545 ? 8'h8f : _GEN_2173; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2175 = 8'h74 == _T_545 ? 8'h92 : _GEN_2174; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2176 = 8'h75 == _T_545 ? 8'h9d : _GEN_2175; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2177 = 8'h76 == _T_545 ? 8'h38 : _GEN_2176; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2178 = 8'h77 == _T_545 ? 8'hf5 : _GEN_2177; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2179 = 8'h78 == _T_545 ? 8'hbc : _GEN_2178; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2180 = 8'h79 == _T_545 ? 8'hb6 : _GEN_2179; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2181 = 8'h7a == _T_545 ? 8'hda : _GEN_2180; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2182 = 8'h7b == _T_545 ? 8'h21 : _GEN_2181; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2183 = 8'h7c == _T_545 ? 8'h10 : _GEN_2182; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2184 = 8'h7d == _T_545 ? 8'hff : _GEN_2183; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2185 = 8'h7e == _T_545 ? 8'hf3 : _GEN_2184; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2186 = 8'h7f == _T_545 ? 8'hd2 : _GEN_2185; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2187 = 8'h80 == _T_545 ? 8'hcd : _GEN_2186; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2188 = 8'h81 == _T_545 ? 8'hc : _GEN_2187; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2189 = 8'h82 == _T_545 ? 8'h13 : _GEN_2188; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2190 = 8'h83 == _T_545 ? 8'hec : _GEN_2189; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2191 = 8'h84 == _T_545 ? 8'h5f : _GEN_2190; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2192 = 8'h85 == _T_545 ? 8'h97 : _GEN_2191; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2193 = 8'h86 == _T_545 ? 8'h44 : _GEN_2192; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2194 = 8'h87 == _T_545 ? 8'h17 : _GEN_2193; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2195 = 8'h88 == _T_545 ? 8'hc4 : _GEN_2194; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2196 = 8'h89 == _T_545 ? 8'ha7 : _GEN_2195; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2197 = 8'h8a == _T_545 ? 8'h7e : _GEN_2196; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2198 = 8'h8b == _T_545 ? 8'h3d : _GEN_2197; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2199 = 8'h8c == _T_545 ? 8'h64 : _GEN_2198; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2200 = 8'h8d == _T_545 ? 8'h5d : _GEN_2199; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2201 = 8'h8e == _T_545 ? 8'h19 : _GEN_2200; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2202 = 8'h8f == _T_545 ? 8'h73 : _GEN_2201; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2203 = 8'h90 == _T_545 ? 8'h60 : _GEN_2202; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2204 = 8'h91 == _T_545 ? 8'h81 : _GEN_2203; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2205 = 8'h92 == _T_545 ? 8'h4f : _GEN_2204; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2206 = 8'h93 == _T_545 ? 8'hdc : _GEN_2205; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2207 = 8'h94 == _T_545 ? 8'h22 : _GEN_2206; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2208 = 8'h95 == _T_545 ? 8'h2a : _GEN_2207; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2209 = 8'h96 == _T_545 ? 8'h90 : _GEN_2208; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2210 = 8'h97 == _T_545 ? 8'h88 : _GEN_2209; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2211 = 8'h98 == _T_545 ? 8'h46 : _GEN_2210; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2212 = 8'h99 == _T_545 ? 8'hee : _GEN_2211; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2213 = 8'h9a == _T_545 ? 8'hb8 : _GEN_2212; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2214 = 8'h9b == _T_545 ? 8'h14 : _GEN_2213; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2215 = 8'h9c == _T_545 ? 8'hde : _GEN_2214; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2216 = 8'h9d == _T_545 ? 8'h5e : _GEN_2215; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2217 = 8'h9e == _T_545 ? 8'hb : _GEN_2216; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2218 = 8'h9f == _T_545 ? 8'hdb : _GEN_2217; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2219 = 8'ha0 == _T_545 ? 8'he0 : _GEN_2218; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2220 = 8'ha1 == _T_545 ? 8'h32 : _GEN_2219; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2221 = 8'ha2 == _T_545 ? 8'h3a : _GEN_2220; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2222 = 8'ha3 == _T_545 ? 8'ha : _GEN_2221; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2223 = 8'ha4 == _T_545 ? 8'h49 : _GEN_2222; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2224 = 8'ha5 == _T_545 ? 8'h6 : _GEN_2223; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2225 = 8'ha6 == _T_545 ? 8'h24 : _GEN_2224; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2226 = 8'ha7 == _T_545 ? 8'h5c : _GEN_2225; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2227 = 8'ha8 == _T_545 ? 8'hc2 : _GEN_2226; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2228 = 8'ha9 == _T_545 ? 8'hd3 : _GEN_2227; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2229 = 8'haa == _T_545 ? 8'hac : _GEN_2228; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2230 = 8'hab == _T_545 ? 8'h62 : _GEN_2229; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2231 = 8'hac == _T_545 ? 8'h91 : _GEN_2230; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2232 = 8'had == _T_545 ? 8'h95 : _GEN_2231; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2233 = 8'hae == _T_545 ? 8'he4 : _GEN_2232; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2234 = 8'haf == _T_545 ? 8'h79 : _GEN_2233; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2235 = 8'hb0 == _T_545 ? 8'he7 : _GEN_2234; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2236 = 8'hb1 == _T_545 ? 8'hc8 : _GEN_2235; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2237 = 8'hb2 == _T_545 ? 8'h37 : _GEN_2236; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2238 = 8'hb3 == _T_545 ? 8'h6d : _GEN_2237; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2239 = 8'hb4 == _T_545 ? 8'h8d : _GEN_2238; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2240 = 8'hb5 == _T_545 ? 8'hd5 : _GEN_2239; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2241 = 8'hb6 == _T_545 ? 8'h4e : _GEN_2240; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2242 = 8'hb7 == _T_545 ? 8'ha9 : _GEN_2241; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2243 = 8'hb8 == _T_545 ? 8'h6c : _GEN_2242; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2244 = 8'hb9 == _T_545 ? 8'h56 : _GEN_2243; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2245 = 8'hba == _T_545 ? 8'hf4 : _GEN_2244; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2246 = 8'hbb == _T_545 ? 8'hea : _GEN_2245; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2247 = 8'hbc == _T_545 ? 8'h65 : _GEN_2246; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2248 = 8'hbd == _T_545 ? 8'h7a : _GEN_2247; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2249 = 8'hbe == _T_545 ? 8'hae : _GEN_2248; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2250 = 8'hbf == _T_545 ? 8'h8 : _GEN_2249; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2251 = 8'hc0 == _T_545 ? 8'hba : _GEN_2250; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2252 = 8'hc1 == _T_545 ? 8'h78 : _GEN_2251; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2253 = 8'hc2 == _T_545 ? 8'h25 : _GEN_2252; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2254 = 8'hc3 == _T_545 ? 8'h2e : _GEN_2253; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2255 = 8'hc4 == _T_545 ? 8'h1c : _GEN_2254; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2256 = 8'hc5 == _T_545 ? 8'ha6 : _GEN_2255; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2257 = 8'hc6 == _T_545 ? 8'hb4 : _GEN_2256; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2258 = 8'hc7 == _T_545 ? 8'hc6 : _GEN_2257; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2259 = 8'hc8 == _T_545 ? 8'he8 : _GEN_2258; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2260 = 8'hc9 == _T_545 ? 8'hdd : _GEN_2259; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2261 = 8'hca == _T_545 ? 8'h74 : _GEN_2260; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2262 = 8'hcb == _T_545 ? 8'h1f : _GEN_2261; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2263 = 8'hcc == _T_545 ? 8'h4b : _GEN_2262; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2264 = 8'hcd == _T_545 ? 8'hbd : _GEN_2263; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2265 = 8'hce == _T_545 ? 8'h8b : _GEN_2264; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2266 = 8'hcf == _T_545 ? 8'h8a : _GEN_2265; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2267 = 8'hd0 == _T_545 ? 8'h70 : _GEN_2266; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2268 = 8'hd1 == _T_545 ? 8'h3e : _GEN_2267; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2269 = 8'hd2 == _T_545 ? 8'hb5 : _GEN_2268; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2270 = 8'hd3 == _T_545 ? 8'h66 : _GEN_2269; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2271 = 8'hd4 == _T_545 ? 8'h48 : _GEN_2270; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2272 = 8'hd5 == _T_545 ? 8'h3 : _GEN_2271; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2273 = 8'hd6 == _T_545 ? 8'hf6 : _GEN_2272; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2274 = 8'hd7 == _T_545 ? 8'he : _GEN_2273; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2275 = 8'hd8 == _T_545 ? 8'h61 : _GEN_2274; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2276 = 8'hd9 == _T_545 ? 8'h35 : _GEN_2275; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2277 = 8'hda == _T_545 ? 8'h57 : _GEN_2276; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2278 = 8'hdb == _T_545 ? 8'hb9 : _GEN_2277; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2279 = 8'hdc == _T_545 ? 8'h86 : _GEN_2278; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2280 = 8'hdd == _T_545 ? 8'hc1 : _GEN_2279; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2281 = 8'hde == _T_545 ? 8'h1d : _GEN_2280; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2282 = 8'hdf == _T_545 ? 8'h9e : _GEN_2281; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2283 = 8'he0 == _T_545 ? 8'he1 : _GEN_2282; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2284 = 8'he1 == _T_545 ? 8'hf8 : _GEN_2283; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2285 = 8'he2 == _T_545 ? 8'h98 : _GEN_2284; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2286 = 8'he3 == _T_545 ? 8'h11 : _GEN_2285; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2287 = 8'he4 == _T_545 ? 8'h69 : _GEN_2286; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2288 = 8'he5 == _T_545 ? 8'hd9 : _GEN_2287; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2289 = 8'he6 == _T_545 ? 8'h8e : _GEN_2288; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2290 = 8'he7 == _T_545 ? 8'h94 : _GEN_2289; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2291 = 8'he8 == _T_545 ? 8'h9b : _GEN_2290; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2292 = 8'he9 == _T_545 ? 8'h1e : _GEN_2291; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2293 = 8'hea == _T_545 ? 8'h87 : _GEN_2292; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2294 = 8'heb == _T_545 ? 8'he9 : _GEN_2293; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2295 = 8'hec == _T_545 ? 8'hce : _GEN_2294; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2296 = 8'hed == _T_545 ? 8'h55 : _GEN_2295; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2297 = 8'hee == _T_545 ? 8'h28 : _GEN_2296; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2298 = 8'hef == _T_545 ? 8'hdf : _GEN_2297; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2299 = 8'hf0 == _T_545 ? 8'h8c : _GEN_2298; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2300 = 8'hf1 == _T_545 ? 8'ha1 : _GEN_2299; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2301 = 8'hf2 == _T_545 ? 8'h89 : _GEN_2300; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2302 = 8'hf3 == _T_545 ? 8'hd : _GEN_2301; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2303 = 8'hf4 == _T_545 ? 8'hbf : _GEN_2302; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2304 = 8'hf5 == _T_545 ? 8'he6 : _GEN_2303; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2305 = 8'hf6 == _T_545 ? 8'h42 : _GEN_2304; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2306 = 8'hf7 == _T_545 ? 8'h68 : _GEN_2305; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2307 = 8'hf8 == _T_545 ? 8'h41 : _GEN_2306; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2308 = 8'hf9 == _T_545 ? 8'h99 : _GEN_2307; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2309 = 8'hfa == _T_545 ? 8'h2d : _GEN_2308; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2310 = 8'hfb == _T_545 ? 8'hf : _GEN_2309; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2311 = 8'hfc == _T_545 ? 8'hb0 : _GEN_2310; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2312 = 8'hfd == _T_545 ? 8'h54 : _GEN_2311; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2313 = 8'hfe == _T_545 ? 8'hbb : _GEN_2312; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2314 = 8'hff == _T_545 ? 8'h16 : _GEN_2313; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2315 = 8'h1 == _T_543 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2316 = 8'h2 == _T_543 ? 8'h77 : _GEN_2315; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2317 = 8'h3 == _T_543 ? 8'h7b : _GEN_2316; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2318 = 8'h4 == _T_543 ? 8'hf2 : _GEN_2317; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2319 = 8'h5 == _T_543 ? 8'h6b : _GEN_2318; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2320 = 8'h6 == _T_543 ? 8'h6f : _GEN_2319; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2321 = 8'h7 == _T_543 ? 8'hc5 : _GEN_2320; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2322 = 8'h8 == _T_543 ? 8'h30 : _GEN_2321; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2323 = 8'h9 == _T_543 ? 8'h1 : _GEN_2322; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2324 = 8'ha == _T_543 ? 8'h67 : _GEN_2323; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2325 = 8'hb == _T_543 ? 8'h2b : _GEN_2324; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2326 = 8'hc == _T_543 ? 8'hfe : _GEN_2325; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2327 = 8'hd == _T_543 ? 8'hd7 : _GEN_2326; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2328 = 8'he == _T_543 ? 8'hab : _GEN_2327; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2329 = 8'hf == _T_543 ? 8'h76 : _GEN_2328; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2330 = 8'h10 == _T_543 ? 8'hca : _GEN_2329; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2331 = 8'h11 == _T_543 ? 8'h82 : _GEN_2330; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2332 = 8'h12 == _T_543 ? 8'hc9 : _GEN_2331; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2333 = 8'h13 == _T_543 ? 8'h7d : _GEN_2332; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2334 = 8'h14 == _T_543 ? 8'hfa : _GEN_2333; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2335 = 8'h15 == _T_543 ? 8'h59 : _GEN_2334; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2336 = 8'h16 == _T_543 ? 8'h47 : _GEN_2335; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2337 = 8'h17 == _T_543 ? 8'hf0 : _GEN_2336; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2338 = 8'h18 == _T_543 ? 8'had : _GEN_2337; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2339 = 8'h19 == _T_543 ? 8'hd4 : _GEN_2338; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2340 = 8'h1a == _T_543 ? 8'ha2 : _GEN_2339; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2341 = 8'h1b == _T_543 ? 8'haf : _GEN_2340; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2342 = 8'h1c == _T_543 ? 8'h9c : _GEN_2341; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2343 = 8'h1d == _T_543 ? 8'ha4 : _GEN_2342; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2344 = 8'h1e == _T_543 ? 8'h72 : _GEN_2343; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2345 = 8'h1f == _T_543 ? 8'hc0 : _GEN_2344; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2346 = 8'h20 == _T_543 ? 8'hb7 : _GEN_2345; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2347 = 8'h21 == _T_543 ? 8'hfd : _GEN_2346; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2348 = 8'h22 == _T_543 ? 8'h93 : _GEN_2347; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2349 = 8'h23 == _T_543 ? 8'h26 : _GEN_2348; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2350 = 8'h24 == _T_543 ? 8'h36 : _GEN_2349; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2351 = 8'h25 == _T_543 ? 8'h3f : _GEN_2350; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2352 = 8'h26 == _T_543 ? 8'hf7 : _GEN_2351; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2353 = 8'h27 == _T_543 ? 8'hcc : _GEN_2352; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2354 = 8'h28 == _T_543 ? 8'h34 : _GEN_2353; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2355 = 8'h29 == _T_543 ? 8'ha5 : _GEN_2354; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2356 = 8'h2a == _T_543 ? 8'he5 : _GEN_2355; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2357 = 8'h2b == _T_543 ? 8'hf1 : _GEN_2356; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2358 = 8'h2c == _T_543 ? 8'h71 : _GEN_2357; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2359 = 8'h2d == _T_543 ? 8'hd8 : _GEN_2358; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2360 = 8'h2e == _T_543 ? 8'h31 : _GEN_2359; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2361 = 8'h2f == _T_543 ? 8'h15 : _GEN_2360; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2362 = 8'h30 == _T_543 ? 8'h4 : _GEN_2361; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2363 = 8'h31 == _T_543 ? 8'hc7 : _GEN_2362; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2364 = 8'h32 == _T_543 ? 8'h23 : _GEN_2363; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2365 = 8'h33 == _T_543 ? 8'hc3 : _GEN_2364; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2366 = 8'h34 == _T_543 ? 8'h18 : _GEN_2365; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2367 = 8'h35 == _T_543 ? 8'h96 : _GEN_2366; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2368 = 8'h36 == _T_543 ? 8'h5 : _GEN_2367; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2369 = 8'h37 == _T_543 ? 8'h9a : _GEN_2368; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2370 = 8'h38 == _T_543 ? 8'h7 : _GEN_2369; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2371 = 8'h39 == _T_543 ? 8'h12 : _GEN_2370; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2372 = 8'h3a == _T_543 ? 8'h80 : _GEN_2371; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2373 = 8'h3b == _T_543 ? 8'he2 : _GEN_2372; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2374 = 8'h3c == _T_543 ? 8'heb : _GEN_2373; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2375 = 8'h3d == _T_543 ? 8'h27 : _GEN_2374; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2376 = 8'h3e == _T_543 ? 8'hb2 : _GEN_2375; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2377 = 8'h3f == _T_543 ? 8'h75 : _GEN_2376; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2378 = 8'h40 == _T_543 ? 8'h9 : _GEN_2377; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2379 = 8'h41 == _T_543 ? 8'h83 : _GEN_2378; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2380 = 8'h42 == _T_543 ? 8'h2c : _GEN_2379; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2381 = 8'h43 == _T_543 ? 8'h1a : _GEN_2380; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2382 = 8'h44 == _T_543 ? 8'h1b : _GEN_2381; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2383 = 8'h45 == _T_543 ? 8'h6e : _GEN_2382; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2384 = 8'h46 == _T_543 ? 8'h5a : _GEN_2383; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2385 = 8'h47 == _T_543 ? 8'ha0 : _GEN_2384; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2386 = 8'h48 == _T_543 ? 8'h52 : _GEN_2385; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2387 = 8'h49 == _T_543 ? 8'h3b : _GEN_2386; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2388 = 8'h4a == _T_543 ? 8'hd6 : _GEN_2387; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2389 = 8'h4b == _T_543 ? 8'hb3 : _GEN_2388; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2390 = 8'h4c == _T_543 ? 8'h29 : _GEN_2389; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2391 = 8'h4d == _T_543 ? 8'he3 : _GEN_2390; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2392 = 8'h4e == _T_543 ? 8'h2f : _GEN_2391; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2393 = 8'h4f == _T_543 ? 8'h84 : _GEN_2392; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2394 = 8'h50 == _T_543 ? 8'h53 : _GEN_2393; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2395 = 8'h51 == _T_543 ? 8'hd1 : _GEN_2394; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2396 = 8'h52 == _T_543 ? 8'h0 : _GEN_2395; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2397 = 8'h53 == _T_543 ? 8'hed : _GEN_2396; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2398 = 8'h54 == _T_543 ? 8'h20 : _GEN_2397; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2399 = 8'h55 == _T_543 ? 8'hfc : _GEN_2398; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2400 = 8'h56 == _T_543 ? 8'hb1 : _GEN_2399; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2401 = 8'h57 == _T_543 ? 8'h5b : _GEN_2400; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2402 = 8'h58 == _T_543 ? 8'h6a : _GEN_2401; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2403 = 8'h59 == _T_543 ? 8'hcb : _GEN_2402; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2404 = 8'h5a == _T_543 ? 8'hbe : _GEN_2403; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2405 = 8'h5b == _T_543 ? 8'h39 : _GEN_2404; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2406 = 8'h5c == _T_543 ? 8'h4a : _GEN_2405; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2407 = 8'h5d == _T_543 ? 8'h4c : _GEN_2406; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2408 = 8'h5e == _T_543 ? 8'h58 : _GEN_2407; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2409 = 8'h5f == _T_543 ? 8'hcf : _GEN_2408; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2410 = 8'h60 == _T_543 ? 8'hd0 : _GEN_2409; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2411 = 8'h61 == _T_543 ? 8'hef : _GEN_2410; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2412 = 8'h62 == _T_543 ? 8'haa : _GEN_2411; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2413 = 8'h63 == _T_543 ? 8'hfb : _GEN_2412; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2414 = 8'h64 == _T_543 ? 8'h43 : _GEN_2413; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2415 = 8'h65 == _T_543 ? 8'h4d : _GEN_2414; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2416 = 8'h66 == _T_543 ? 8'h33 : _GEN_2415; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2417 = 8'h67 == _T_543 ? 8'h85 : _GEN_2416; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2418 = 8'h68 == _T_543 ? 8'h45 : _GEN_2417; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2419 = 8'h69 == _T_543 ? 8'hf9 : _GEN_2418; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2420 = 8'h6a == _T_543 ? 8'h2 : _GEN_2419; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2421 = 8'h6b == _T_543 ? 8'h7f : _GEN_2420; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2422 = 8'h6c == _T_543 ? 8'h50 : _GEN_2421; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2423 = 8'h6d == _T_543 ? 8'h3c : _GEN_2422; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2424 = 8'h6e == _T_543 ? 8'h9f : _GEN_2423; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2425 = 8'h6f == _T_543 ? 8'ha8 : _GEN_2424; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2426 = 8'h70 == _T_543 ? 8'h51 : _GEN_2425; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2427 = 8'h71 == _T_543 ? 8'ha3 : _GEN_2426; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2428 = 8'h72 == _T_543 ? 8'h40 : _GEN_2427; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2429 = 8'h73 == _T_543 ? 8'h8f : _GEN_2428; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2430 = 8'h74 == _T_543 ? 8'h92 : _GEN_2429; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2431 = 8'h75 == _T_543 ? 8'h9d : _GEN_2430; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2432 = 8'h76 == _T_543 ? 8'h38 : _GEN_2431; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2433 = 8'h77 == _T_543 ? 8'hf5 : _GEN_2432; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2434 = 8'h78 == _T_543 ? 8'hbc : _GEN_2433; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2435 = 8'h79 == _T_543 ? 8'hb6 : _GEN_2434; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2436 = 8'h7a == _T_543 ? 8'hda : _GEN_2435; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2437 = 8'h7b == _T_543 ? 8'h21 : _GEN_2436; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2438 = 8'h7c == _T_543 ? 8'h10 : _GEN_2437; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2439 = 8'h7d == _T_543 ? 8'hff : _GEN_2438; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2440 = 8'h7e == _T_543 ? 8'hf3 : _GEN_2439; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2441 = 8'h7f == _T_543 ? 8'hd2 : _GEN_2440; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2442 = 8'h80 == _T_543 ? 8'hcd : _GEN_2441; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2443 = 8'h81 == _T_543 ? 8'hc : _GEN_2442; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2444 = 8'h82 == _T_543 ? 8'h13 : _GEN_2443; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2445 = 8'h83 == _T_543 ? 8'hec : _GEN_2444; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2446 = 8'h84 == _T_543 ? 8'h5f : _GEN_2445; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2447 = 8'h85 == _T_543 ? 8'h97 : _GEN_2446; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2448 = 8'h86 == _T_543 ? 8'h44 : _GEN_2447; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2449 = 8'h87 == _T_543 ? 8'h17 : _GEN_2448; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2450 = 8'h88 == _T_543 ? 8'hc4 : _GEN_2449; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2451 = 8'h89 == _T_543 ? 8'ha7 : _GEN_2450; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2452 = 8'h8a == _T_543 ? 8'h7e : _GEN_2451; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2453 = 8'h8b == _T_543 ? 8'h3d : _GEN_2452; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2454 = 8'h8c == _T_543 ? 8'h64 : _GEN_2453; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2455 = 8'h8d == _T_543 ? 8'h5d : _GEN_2454; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2456 = 8'h8e == _T_543 ? 8'h19 : _GEN_2455; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2457 = 8'h8f == _T_543 ? 8'h73 : _GEN_2456; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2458 = 8'h90 == _T_543 ? 8'h60 : _GEN_2457; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2459 = 8'h91 == _T_543 ? 8'h81 : _GEN_2458; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2460 = 8'h92 == _T_543 ? 8'h4f : _GEN_2459; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2461 = 8'h93 == _T_543 ? 8'hdc : _GEN_2460; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2462 = 8'h94 == _T_543 ? 8'h22 : _GEN_2461; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2463 = 8'h95 == _T_543 ? 8'h2a : _GEN_2462; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2464 = 8'h96 == _T_543 ? 8'h90 : _GEN_2463; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2465 = 8'h97 == _T_543 ? 8'h88 : _GEN_2464; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2466 = 8'h98 == _T_543 ? 8'h46 : _GEN_2465; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2467 = 8'h99 == _T_543 ? 8'hee : _GEN_2466; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2468 = 8'h9a == _T_543 ? 8'hb8 : _GEN_2467; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2469 = 8'h9b == _T_543 ? 8'h14 : _GEN_2468; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2470 = 8'h9c == _T_543 ? 8'hde : _GEN_2469; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2471 = 8'h9d == _T_543 ? 8'h5e : _GEN_2470; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2472 = 8'h9e == _T_543 ? 8'hb : _GEN_2471; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2473 = 8'h9f == _T_543 ? 8'hdb : _GEN_2472; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2474 = 8'ha0 == _T_543 ? 8'he0 : _GEN_2473; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2475 = 8'ha1 == _T_543 ? 8'h32 : _GEN_2474; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2476 = 8'ha2 == _T_543 ? 8'h3a : _GEN_2475; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2477 = 8'ha3 == _T_543 ? 8'ha : _GEN_2476; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2478 = 8'ha4 == _T_543 ? 8'h49 : _GEN_2477; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2479 = 8'ha5 == _T_543 ? 8'h6 : _GEN_2478; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2480 = 8'ha6 == _T_543 ? 8'h24 : _GEN_2479; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2481 = 8'ha7 == _T_543 ? 8'h5c : _GEN_2480; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2482 = 8'ha8 == _T_543 ? 8'hc2 : _GEN_2481; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2483 = 8'ha9 == _T_543 ? 8'hd3 : _GEN_2482; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2484 = 8'haa == _T_543 ? 8'hac : _GEN_2483; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2485 = 8'hab == _T_543 ? 8'h62 : _GEN_2484; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2486 = 8'hac == _T_543 ? 8'h91 : _GEN_2485; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2487 = 8'had == _T_543 ? 8'h95 : _GEN_2486; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2488 = 8'hae == _T_543 ? 8'he4 : _GEN_2487; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2489 = 8'haf == _T_543 ? 8'h79 : _GEN_2488; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2490 = 8'hb0 == _T_543 ? 8'he7 : _GEN_2489; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2491 = 8'hb1 == _T_543 ? 8'hc8 : _GEN_2490; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2492 = 8'hb2 == _T_543 ? 8'h37 : _GEN_2491; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2493 = 8'hb3 == _T_543 ? 8'h6d : _GEN_2492; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2494 = 8'hb4 == _T_543 ? 8'h8d : _GEN_2493; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2495 = 8'hb5 == _T_543 ? 8'hd5 : _GEN_2494; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2496 = 8'hb6 == _T_543 ? 8'h4e : _GEN_2495; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2497 = 8'hb7 == _T_543 ? 8'ha9 : _GEN_2496; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2498 = 8'hb8 == _T_543 ? 8'h6c : _GEN_2497; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2499 = 8'hb9 == _T_543 ? 8'h56 : _GEN_2498; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2500 = 8'hba == _T_543 ? 8'hf4 : _GEN_2499; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2501 = 8'hbb == _T_543 ? 8'hea : _GEN_2500; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2502 = 8'hbc == _T_543 ? 8'h65 : _GEN_2501; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2503 = 8'hbd == _T_543 ? 8'h7a : _GEN_2502; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2504 = 8'hbe == _T_543 ? 8'hae : _GEN_2503; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2505 = 8'hbf == _T_543 ? 8'h8 : _GEN_2504; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2506 = 8'hc0 == _T_543 ? 8'hba : _GEN_2505; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2507 = 8'hc1 == _T_543 ? 8'h78 : _GEN_2506; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2508 = 8'hc2 == _T_543 ? 8'h25 : _GEN_2507; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2509 = 8'hc3 == _T_543 ? 8'h2e : _GEN_2508; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2510 = 8'hc4 == _T_543 ? 8'h1c : _GEN_2509; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2511 = 8'hc5 == _T_543 ? 8'ha6 : _GEN_2510; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2512 = 8'hc6 == _T_543 ? 8'hb4 : _GEN_2511; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2513 = 8'hc7 == _T_543 ? 8'hc6 : _GEN_2512; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2514 = 8'hc8 == _T_543 ? 8'he8 : _GEN_2513; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2515 = 8'hc9 == _T_543 ? 8'hdd : _GEN_2514; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2516 = 8'hca == _T_543 ? 8'h74 : _GEN_2515; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2517 = 8'hcb == _T_543 ? 8'h1f : _GEN_2516; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2518 = 8'hcc == _T_543 ? 8'h4b : _GEN_2517; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2519 = 8'hcd == _T_543 ? 8'hbd : _GEN_2518; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2520 = 8'hce == _T_543 ? 8'h8b : _GEN_2519; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2521 = 8'hcf == _T_543 ? 8'h8a : _GEN_2520; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2522 = 8'hd0 == _T_543 ? 8'h70 : _GEN_2521; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2523 = 8'hd1 == _T_543 ? 8'h3e : _GEN_2522; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2524 = 8'hd2 == _T_543 ? 8'hb5 : _GEN_2523; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2525 = 8'hd3 == _T_543 ? 8'h66 : _GEN_2524; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2526 = 8'hd4 == _T_543 ? 8'h48 : _GEN_2525; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2527 = 8'hd5 == _T_543 ? 8'h3 : _GEN_2526; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2528 = 8'hd6 == _T_543 ? 8'hf6 : _GEN_2527; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2529 = 8'hd7 == _T_543 ? 8'he : _GEN_2528; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2530 = 8'hd8 == _T_543 ? 8'h61 : _GEN_2529; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2531 = 8'hd9 == _T_543 ? 8'h35 : _GEN_2530; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2532 = 8'hda == _T_543 ? 8'h57 : _GEN_2531; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2533 = 8'hdb == _T_543 ? 8'hb9 : _GEN_2532; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2534 = 8'hdc == _T_543 ? 8'h86 : _GEN_2533; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2535 = 8'hdd == _T_543 ? 8'hc1 : _GEN_2534; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2536 = 8'hde == _T_543 ? 8'h1d : _GEN_2535; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2537 = 8'hdf == _T_543 ? 8'h9e : _GEN_2536; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2538 = 8'he0 == _T_543 ? 8'he1 : _GEN_2537; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2539 = 8'he1 == _T_543 ? 8'hf8 : _GEN_2538; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2540 = 8'he2 == _T_543 ? 8'h98 : _GEN_2539; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2541 = 8'he3 == _T_543 ? 8'h11 : _GEN_2540; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2542 = 8'he4 == _T_543 ? 8'h69 : _GEN_2541; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2543 = 8'he5 == _T_543 ? 8'hd9 : _GEN_2542; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2544 = 8'he6 == _T_543 ? 8'h8e : _GEN_2543; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2545 = 8'he7 == _T_543 ? 8'h94 : _GEN_2544; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2546 = 8'he8 == _T_543 ? 8'h9b : _GEN_2545; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2547 = 8'he9 == _T_543 ? 8'h1e : _GEN_2546; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2548 = 8'hea == _T_543 ? 8'h87 : _GEN_2547; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2549 = 8'heb == _T_543 ? 8'he9 : _GEN_2548; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2550 = 8'hec == _T_543 ? 8'hce : _GEN_2549; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2551 = 8'hed == _T_543 ? 8'h55 : _GEN_2550; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2552 = 8'hee == _T_543 ? 8'h28 : _GEN_2551; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2553 = 8'hef == _T_543 ? 8'hdf : _GEN_2552; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2554 = 8'hf0 == _T_543 ? 8'h8c : _GEN_2553; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2555 = 8'hf1 == _T_543 ? 8'ha1 : _GEN_2554; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2556 = 8'hf2 == _T_543 ? 8'h89 : _GEN_2555; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2557 = 8'hf3 == _T_543 ? 8'hd : _GEN_2556; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2558 = 8'hf4 == _T_543 ? 8'hbf : _GEN_2557; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2559 = 8'hf5 == _T_543 ? 8'he6 : _GEN_2558; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2560 = 8'hf6 == _T_543 ? 8'h42 : _GEN_2559; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2561 = 8'hf7 == _T_543 ? 8'h68 : _GEN_2560; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2562 = 8'hf8 == _T_543 ? 8'h41 : _GEN_2561; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2563 = 8'hf9 == _T_543 ? 8'h99 : _GEN_2562; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2564 = 8'hfa == _T_543 ? 8'h2d : _GEN_2563; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2565 = 8'hfb == _T_543 ? 8'hf : _GEN_2564; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2566 = 8'hfc == _T_543 ? 8'hb0 : _GEN_2565; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2567 = 8'hfd == _T_543 ? 8'h54 : _GEN_2566; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2568 = 8'hfe == _T_543 ? 8'hbb : _GEN_2567; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2569 = 8'hff == _T_543 ? 8'h16 : _GEN_2568; // @[Cat.scala 30:58:@2080.4]
  assign _T_551 = {_GEN_2314,_GEN_2569}; // @[Cat.scala 30:58:@2080.4]
  assign _GEN_2570 = 8'h1 == _T_549 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2571 = 8'h2 == _T_549 ? 8'h77 : _GEN_2570; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2572 = 8'h3 == _T_549 ? 8'h7b : _GEN_2571; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2573 = 8'h4 == _T_549 ? 8'hf2 : _GEN_2572; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2574 = 8'h5 == _T_549 ? 8'h6b : _GEN_2573; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2575 = 8'h6 == _T_549 ? 8'h6f : _GEN_2574; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2576 = 8'h7 == _T_549 ? 8'hc5 : _GEN_2575; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2577 = 8'h8 == _T_549 ? 8'h30 : _GEN_2576; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2578 = 8'h9 == _T_549 ? 8'h1 : _GEN_2577; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2579 = 8'ha == _T_549 ? 8'h67 : _GEN_2578; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2580 = 8'hb == _T_549 ? 8'h2b : _GEN_2579; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2581 = 8'hc == _T_549 ? 8'hfe : _GEN_2580; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2582 = 8'hd == _T_549 ? 8'hd7 : _GEN_2581; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2583 = 8'he == _T_549 ? 8'hab : _GEN_2582; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2584 = 8'hf == _T_549 ? 8'h76 : _GEN_2583; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2585 = 8'h10 == _T_549 ? 8'hca : _GEN_2584; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2586 = 8'h11 == _T_549 ? 8'h82 : _GEN_2585; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2587 = 8'h12 == _T_549 ? 8'hc9 : _GEN_2586; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2588 = 8'h13 == _T_549 ? 8'h7d : _GEN_2587; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2589 = 8'h14 == _T_549 ? 8'hfa : _GEN_2588; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2590 = 8'h15 == _T_549 ? 8'h59 : _GEN_2589; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2591 = 8'h16 == _T_549 ? 8'h47 : _GEN_2590; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2592 = 8'h17 == _T_549 ? 8'hf0 : _GEN_2591; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2593 = 8'h18 == _T_549 ? 8'had : _GEN_2592; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2594 = 8'h19 == _T_549 ? 8'hd4 : _GEN_2593; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2595 = 8'h1a == _T_549 ? 8'ha2 : _GEN_2594; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2596 = 8'h1b == _T_549 ? 8'haf : _GEN_2595; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2597 = 8'h1c == _T_549 ? 8'h9c : _GEN_2596; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2598 = 8'h1d == _T_549 ? 8'ha4 : _GEN_2597; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2599 = 8'h1e == _T_549 ? 8'h72 : _GEN_2598; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2600 = 8'h1f == _T_549 ? 8'hc0 : _GEN_2599; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2601 = 8'h20 == _T_549 ? 8'hb7 : _GEN_2600; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2602 = 8'h21 == _T_549 ? 8'hfd : _GEN_2601; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2603 = 8'h22 == _T_549 ? 8'h93 : _GEN_2602; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2604 = 8'h23 == _T_549 ? 8'h26 : _GEN_2603; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2605 = 8'h24 == _T_549 ? 8'h36 : _GEN_2604; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2606 = 8'h25 == _T_549 ? 8'h3f : _GEN_2605; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2607 = 8'h26 == _T_549 ? 8'hf7 : _GEN_2606; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2608 = 8'h27 == _T_549 ? 8'hcc : _GEN_2607; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2609 = 8'h28 == _T_549 ? 8'h34 : _GEN_2608; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2610 = 8'h29 == _T_549 ? 8'ha5 : _GEN_2609; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2611 = 8'h2a == _T_549 ? 8'he5 : _GEN_2610; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2612 = 8'h2b == _T_549 ? 8'hf1 : _GEN_2611; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2613 = 8'h2c == _T_549 ? 8'h71 : _GEN_2612; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2614 = 8'h2d == _T_549 ? 8'hd8 : _GEN_2613; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2615 = 8'h2e == _T_549 ? 8'h31 : _GEN_2614; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2616 = 8'h2f == _T_549 ? 8'h15 : _GEN_2615; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2617 = 8'h30 == _T_549 ? 8'h4 : _GEN_2616; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2618 = 8'h31 == _T_549 ? 8'hc7 : _GEN_2617; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2619 = 8'h32 == _T_549 ? 8'h23 : _GEN_2618; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2620 = 8'h33 == _T_549 ? 8'hc3 : _GEN_2619; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2621 = 8'h34 == _T_549 ? 8'h18 : _GEN_2620; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2622 = 8'h35 == _T_549 ? 8'h96 : _GEN_2621; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2623 = 8'h36 == _T_549 ? 8'h5 : _GEN_2622; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2624 = 8'h37 == _T_549 ? 8'h9a : _GEN_2623; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2625 = 8'h38 == _T_549 ? 8'h7 : _GEN_2624; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2626 = 8'h39 == _T_549 ? 8'h12 : _GEN_2625; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2627 = 8'h3a == _T_549 ? 8'h80 : _GEN_2626; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2628 = 8'h3b == _T_549 ? 8'he2 : _GEN_2627; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2629 = 8'h3c == _T_549 ? 8'heb : _GEN_2628; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2630 = 8'h3d == _T_549 ? 8'h27 : _GEN_2629; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2631 = 8'h3e == _T_549 ? 8'hb2 : _GEN_2630; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2632 = 8'h3f == _T_549 ? 8'h75 : _GEN_2631; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2633 = 8'h40 == _T_549 ? 8'h9 : _GEN_2632; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2634 = 8'h41 == _T_549 ? 8'h83 : _GEN_2633; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2635 = 8'h42 == _T_549 ? 8'h2c : _GEN_2634; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2636 = 8'h43 == _T_549 ? 8'h1a : _GEN_2635; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2637 = 8'h44 == _T_549 ? 8'h1b : _GEN_2636; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2638 = 8'h45 == _T_549 ? 8'h6e : _GEN_2637; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2639 = 8'h46 == _T_549 ? 8'h5a : _GEN_2638; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2640 = 8'h47 == _T_549 ? 8'ha0 : _GEN_2639; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2641 = 8'h48 == _T_549 ? 8'h52 : _GEN_2640; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2642 = 8'h49 == _T_549 ? 8'h3b : _GEN_2641; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2643 = 8'h4a == _T_549 ? 8'hd6 : _GEN_2642; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2644 = 8'h4b == _T_549 ? 8'hb3 : _GEN_2643; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2645 = 8'h4c == _T_549 ? 8'h29 : _GEN_2644; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2646 = 8'h4d == _T_549 ? 8'he3 : _GEN_2645; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2647 = 8'h4e == _T_549 ? 8'h2f : _GEN_2646; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2648 = 8'h4f == _T_549 ? 8'h84 : _GEN_2647; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2649 = 8'h50 == _T_549 ? 8'h53 : _GEN_2648; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2650 = 8'h51 == _T_549 ? 8'hd1 : _GEN_2649; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2651 = 8'h52 == _T_549 ? 8'h0 : _GEN_2650; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2652 = 8'h53 == _T_549 ? 8'hed : _GEN_2651; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2653 = 8'h54 == _T_549 ? 8'h20 : _GEN_2652; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2654 = 8'h55 == _T_549 ? 8'hfc : _GEN_2653; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2655 = 8'h56 == _T_549 ? 8'hb1 : _GEN_2654; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2656 = 8'h57 == _T_549 ? 8'h5b : _GEN_2655; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2657 = 8'h58 == _T_549 ? 8'h6a : _GEN_2656; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2658 = 8'h59 == _T_549 ? 8'hcb : _GEN_2657; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2659 = 8'h5a == _T_549 ? 8'hbe : _GEN_2658; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2660 = 8'h5b == _T_549 ? 8'h39 : _GEN_2659; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2661 = 8'h5c == _T_549 ? 8'h4a : _GEN_2660; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2662 = 8'h5d == _T_549 ? 8'h4c : _GEN_2661; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2663 = 8'h5e == _T_549 ? 8'h58 : _GEN_2662; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2664 = 8'h5f == _T_549 ? 8'hcf : _GEN_2663; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2665 = 8'h60 == _T_549 ? 8'hd0 : _GEN_2664; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2666 = 8'h61 == _T_549 ? 8'hef : _GEN_2665; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2667 = 8'h62 == _T_549 ? 8'haa : _GEN_2666; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2668 = 8'h63 == _T_549 ? 8'hfb : _GEN_2667; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2669 = 8'h64 == _T_549 ? 8'h43 : _GEN_2668; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2670 = 8'h65 == _T_549 ? 8'h4d : _GEN_2669; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2671 = 8'h66 == _T_549 ? 8'h33 : _GEN_2670; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2672 = 8'h67 == _T_549 ? 8'h85 : _GEN_2671; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2673 = 8'h68 == _T_549 ? 8'h45 : _GEN_2672; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2674 = 8'h69 == _T_549 ? 8'hf9 : _GEN_2673; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2675 = 8'h6a == _T_549 ? 8'h2 : _GEN_2674; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2676 = 8'h6b == _T_549 ? 8'h7f : _GEN_2675; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2677 = 8'h6c == _T_549 ? 8'h50 : _GEN_2676; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2678 = 8'h6d == _T_549 ? 8'h3c : _GEN_2677; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2679 = 8'h6e == _T_549 ? 8'h9f : _GEN_2678; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2680 = 8'h6f == _T_549 ? 8'ha8 : _GEN_2679; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2681 = 8'h70 == _T_549 ? 8'h51 : _GEN_2680; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2682 = 8'h71 == _T_549 ? 8'ha3 : _GEN_2681; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2683 = 8'h72 == _T_549 ? 8'h40 : _GEN_2682; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2684 = 8'h73 == _T_549 ? 8'h8f : _GEN_2683; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2685 = 8'h74 == _T_549 ? 8'h92 : _GEN_2684; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2686 = 8'h75 == _T_549 ? 8'h9d : _GEN_2685; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2687 = 8'h76 == _T_549 ? 8'h38 : _GEN_2686; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2688 = 8'h77 == _T_549 ? 8'hf5 : _GEN_2687; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2689 = 8'h78 == _T_549 ? 8'hbc : _GEN_2688; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2690 = 8'h79 == _T_549 ? 8'hb6 : _GEN_2689; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2691 = 8'h7a == _T_549 ? 8'hda : _GEN_2690; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2692 = 8'h7b == _T_549 ? 8'h21 : _GEN_2691; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2693 = 8'h7c == _T_549 ? 8'h10 : _GEN_2692; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2694 = 8'h7d == _T_549 ? 8'hff : _GEN_2693; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2695 = 8'h7e == _T_549 ? 8'hf3 : _GEN_2694; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2696 = 8'h7f == _T_549 ? 8'hd2 : _GEN_2695; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2697 = 8'h80 == _T_549 ? 8'hcd : _GEN_2696; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2698 = 8'h81 == _T_549 ? 8'hc : _GEN_2697; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2699 = 8'h82 == _T_549 ? 8'h13 : _GEN_2698; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2700 = 8'h83 == _T_549 ? 8'hec : _GEN_2699; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2701 = 8'h84 == _T_549 ? 8'h5f : _GEN_2700; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2702 = 8'h85 == _T_549 ? 8'h97 : _GEN_2701; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2703 = 8'h86 == _T_549 ? 8'h44 : _GEN_2702; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2704 = 8'h87 == _T_549 ? 8'h17 : _GEN_2703; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2705 = 8'h88 == _T_549 ? 8'hc4 : _GEN_2704; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2706 = 8'h89 == _T_549 ? 8'ha7 : _GEN_2705; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2707 = 8'h8a == _T_549 ? 8'h7e : _GEN_2706; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2708 = 8'h8b == _T_549 ? 8'h3d : _GEN_2707; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2709 = 8'h8c == _T_549 ? 8'h64 : _GEN_2708; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2710 = 8'h8d == _T_549 ? 8'h5d : _GEN_2709; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2711 = 8'h8e == _T_549 ? 8'h19 : _GEN_2710; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2712 = 8'h8f == _T_549 ? 8'h73 : _GEN_2711; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2713 = 8'h90 == _T_549 ? 8'h60 : _GEN_2712; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2714 = 8'h91 == _T_549 ? 8'h81 : _GEN_2713; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2715 = 8'h92 == _T_549 ? 8'h4f : _GEN_2714; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2716 = 8'h93 == _T_549 ? 8'hdc : _GEN_2715; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2717 = 8'h94 == _T_549 ? 8'h22 : _GEN_2716; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2718 = 8'h95 == _T_549 ? 8'h2a : _GEN_2717; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2719 = 8'h96 == _T_549 ? 8'h90 : _GEN_2718; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2720 = 8'h97 == _T_549 ? 8'h88 : _GEN_2719; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2721 = 8'h98 == _T_549 ? 8'h46 : _GEN_2720; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2722 = 8'h99 == _T_549 ? 8'hee : _GEN_2721; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2723 = 8'h9a == _T_549 ? 8'hb8 : _GEN_2722; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2724 = 8'h9b == _T_549 ? 8'h14 : _GEN_2723; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2725 = 8'h9c == _T_549 ? 8'hde : _GEN_2724; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2726 = 8'h9d == _T_549 ? 8'h5e : _GEN_2725; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2727 = 8'h9e == _T_549 ? 8'hb : _GEN_2726; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2728 = 8'h9f == _T_549 ? 8'hdb : _GEN_2727; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2729 = 8'ha0 == _T_549 ? 8'he0 : _GEN_2728; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2730 = 8'ha1 == _T_549 ? 8'h32 : _GEN_2729; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2731 = 8'ha2 == _T_549 ? 8'h3a : _GEN_2730; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2732 = 8'ha3 == _T_549 ? 8'ha : _GEN_2731; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2733 = 8'ha4 == _T_549 ? 8'h49 : _GEN_2732; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2734 = 8'ha5 == _T_549 ? 8'h6 : _GEN_2733; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2735 = 8'ha6 == _T_549 ? 8'h24 : _GEN_2734; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2736 = 8'ha7 == _T_549 ? 8'h5c : _GEN_2735; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2737 = 8'ha8 == _T_549 ? 8'hc2 : _GEN_2736; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2738 = 8'ha9 == _T_549 ? 8'hd3 : _GEN_2737; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2739 = 8'haa == _T_549 ? 8'hac : _GEN_2738; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2740 = 8'hab == _T_549 ? 8'h62 : _GEN_2739; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2741 = 8'hac == _T_549 ? 8'h91 : _GEN_2740; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2742 = 8'had == _T_549 ? 8'h95 : _GEN_2741; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2743 = 8'hae == _T_549 ? 8'he4 : _GEN_2742; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2744 = 8'haf == _T_549 ? 8'h79 : _GEN_2743; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2745 = 8'hb0 == _T_549 ? 8'he7 : _GEN_2744; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2746 = 8'hb1 == _T_549 ? 8'hc8 : _GEN_2745; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2747 = 8'hb2 == _T_549 ? 8'h37 : _GEN_2746; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2748 = 8'hb3 == _T_549 ? 8'h6d : _GEN_2747; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2749 = 8'hb4 == _T_549 ? 8'h8d : _GEN_2748; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2750 = 8'hb5 == _T_549 ? 8'hd5 : _GEN_2749; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2751 = 8'hb6 == _T_549 ? 8'h4e : _GEN_2750; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2752 = 8'hb7 == _T_549 ? 8'ha9 : _GEN_2751; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2753 = 8'hb8 == _T_549 ? 8'h6c : _GEN_2752; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2754 = 8'hb9 == _T_549 ? 8'h56 : _GEN_2753; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2755 = 8'hba == _T_549 ? 8'hf4 : _GEN_2754; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2756 = 8'hbb == _T_549 ? 8'hea : _GEN_2755; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2757 = 8'hbc == _T_549 ? 8'h65 : _GEN_2756; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2758 = 8'hbd == _T_549 ? 8'h7a : _GEN_2757; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2759 = 8'hbe == _T_549 ? 8'hae : _GEN_2758; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2760 = 8'hbf == _T_549 ? 8'h8 : _GEN_2759; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2761 = 8'hc0 == _T_549 ? 8'hba : _GEN_2760; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2762 = 8'hc1 == _T_549 ? 8'h78 : _GEN_2761; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2763 = 8'hc2 == _T_549 ? 8'h25 : _GEN_2762; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2764 = 8'hc3 == _T_549 ? 8'h2e : _GEN_2763; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2765 = 8'hc4 == _T_549 ? 8'h1c : _GEN_2764; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2766 = 8'hc5 == _T_549 ? 8'ha6 : _GEN_2765; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2767 = 8'hc6 == _T_549 ? 8'hb4 : _GEN_2766; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2768 = 8'hc7 == _T_549 ? 8'hc6 : _GEN_2767; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2769 = 8'hc8 == _T_549 ? 8'he8 : _GEN_2768; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2770 = 8'hc9 == _T_549 ? 8'hdd : _GEN_2769; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2771 = 8'hca == _T_549 ? 8'h74 : _GEN_2770; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2772 = 8'hcb == _T_549 ? 8'h1f : _GEN_2771; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2773 = 8'hcc == _T_549 ? 8'h4b : _GEN_2772; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2774 = 8'hcd == _T_549 ? 8'hbd : _GEN_2773; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2775 = 8'hce == _T_549 ? 8'h8b : _GEN_2774; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2776 = 8'hcf == _T_549 ? 8'h8a : _GEN_2775; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2777 = 8'hd0 == _T_549 ? 8'h70 : _GEN_2776; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2778 = 8'hd1 == _T_549 ? 8'h3e : _GEN_2777; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2779 = 8'hd2 == _T_549 ? 8'hb5 : _GEN_2778; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2780 = 8'hd3 == _T_549 ? 8'h66 : _GEN_2779; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2781 = 8'hd4 == _T_549 ? 8'h48 : _GEN_2780; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2782 = 8'hd5 == _T_549 ? 8'h3 : _GEN_2781; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2783 = 8'hd6 == _T_549 ? 8'hf6 : _GEN_2782; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2784 = 8'hd7 == _T_549 ? 8'he : _GEN_2783; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2785 = 8'hd8 == _T_549 ? 8'h61 : _GEN_2784; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2786 = 8'hd9 == _T_549 ? 8'h35 : _GEN_2785; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2787 = 8'hda == _T_549 ? 8'h57 : _GEN_2786; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2788 = 8'hdb == _T_549 ? 8'hb9 : _GEN_2787; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2789 = 8'hdc == _T_549 ? 8'h86 : _GEN_2788; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2790 = 8'hdd == _T_549 ? 8'hc1 : _GEN_2789; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2791 = 8'hde == _T_549 ? 8'h1d : _GEN_2790; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2792 = 8'hdf == _T_549 ? 8'h9e : _GEN_2791; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2793 = 8'he0 == _T_549 ? 8'he1 : _GEN_2792; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2794 = 8'he1 == _T_549 ? 8'hf8 : _GEN_2793; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2795 = 8'he2 == _T_549 ? 8'h98 : _GEN_2794; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2796 = 8'he3 == _T_549 ? 8'h11 : _GEN_2795; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2797 = 8'he4 == _T_549 ? 8'h69 : _GEN_2796; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2798 = 8'he5 == _T_549 ? 8'hd9 : _GEN_2797; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2799 = 8'he6 == _T_549 ? 8'h8e : _GEN_2798; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2800 = 8'he7 == _T_549 ? 8'h94 : _GEN_2799; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2801 = 8'he8 == _T_549 ? 8'h9b : _GEN_2800; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2802 = 8'he9 == _T_549 ? 8'h1e : _GEN_2801; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2803 = 8'hea == _T_549 ? 8'h87 : _GEN_2802; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2804 = 8'heb == _T_549 ? 8'he9 : _GEN_2803; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2805 = 8'hec == _T_549 ? 8'hce : _GEN_2804; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2806 = 8'hed == _T_549 ? 8'h55 : _GEN_2805; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2807 = 8'hee == _T_549 ? 8'h28 : _GEN_2806; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2808 = 8'hef == _T_549 ? 8'hdf : _GEN_2807; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2809 = 8'hf0 == _T_549 ? 8'h8c : _GEN_2808; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2810 = 8'hf1 == _T_549 ? 8'ha1 : _GEN_2809; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2811 = 8'hf2 == _T_549 ? 8'h89 : _GEN_2810; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2812 = 8'hf3 == _T_549 ? 8'hd : _GEN_2811; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2813 = 8'hf4 == _T_549 ? 8'hbf : _GEN_2812; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2814 = 8'hf5 == _T_549 ? 8'he6 : _GEN_2813; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2815 = 8'hf6 == _T_549 ? 8'h42 : _GEN_2814; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2816 = 8'hf7 == _T_549 ? 8'h68 : _GEN_2815; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2817 = 8'hf8 == _T_549 ? 8'h41 : _GEN_2816; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2818 = 8'hf9 == _T_549 ? 8'h99 : _GEN_2817; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2819 = 8'hfa == _T_549 ? 8'h2d : _GEN_2818; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2820 = 8'hfb == _T_549 ? 8'hf : _GEN_2819; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2821 = 8'hfc == _T_549 ? 8'hb0 : _GEN_2820; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2822 = 8'hfd == _T_549 ? 8'h54 : _GEN_2821; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2823 = 8'hfe == _T_549 ? 8'hbb : _GEN_2822; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2824 = 8'hff == _T_549 ? 8'h16 : _GEN_2823; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2825 = 8'h1 == _T_547 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2826 = 8'h2 == _T_547 ? 8'h77 : _GEN_2825; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2827 = 8'h3 == _T_547 ? 8'h7b : _GEN_2826; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2828 = 8'h4 == _T_547 ? 8'hf2 : _GEN_2827; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2829 = 8'h5 == _T_547 ? 8'h6b : _GEN_2828; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2830 = 8'h6 == _T_547 ? 8'h6f : _GEN_2829; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2831 = 8'h7 == _T_547 ? 8'hc5 : _GEN_2830; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2832 = 8'h8 == _T_547 ? 8'h30 : _GEN_2831; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2833 = 8'h9 == _T_547 ? 8'h1 : _GEN_2832; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2834 = 8'ha == _T_547 ? 8'h67 : _GEN_2833; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2835 = 8'hb == _T_547 ? 8'h2b : _GEN_2834; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2836 = 8'hc == _T_547 ? 8'hfe : _GEN_2835; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2837 = 8'hd == _T_547 ? 8'hd7 : _GEN_2836; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2838 = 8'he == _T_547 ? 8'hab : _GEN_2837; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2839 = 8'hf == _T_547 ? 8'h76 : _GEN_2838; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2840 = 8'h10 == _T_547 ? 8'hca : _GEN_2839; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2841 = 8'h11 == _T_547 ? 8'h82 : _GEN_2840; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2842 = 8'h12 == _T_547 ? 8'hc9 : _GEN_2841; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2843 = 8'h13 == _T_547 ? 8'h7d : _GEN_2842; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2844 = 8'h14 == _T_547 ? 8'hfa : _GEN_2843; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2845 = 8'h15 == _T_547 ? 8'h59 : _GEN_2844; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2846 = 8'h16 == _T_547 ? 8'h47 : _GEN_2845; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2847 = 8'h17 == _T_547 ? 8'hf0 : _GEN_2846; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2848 = 8'h18 == _T_547 ? 8'had : _GEN_2847; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2849 = 8'h19 == _T_547 ? 8'hd4 : _GEN_2848; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2850 = 8'h1a == _T_547 ? 8'ha2 : _GEN_2849; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2851 = 8'h1b == _T_547 ? 8'haf : _GEN_2850; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2852 = 8'h1c == _T_547 ? 8'h9c : _GEN_2851; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2853 = 8'h1d == _T_547 ? 8'ha4 : _GEN_2852; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2854 = 8'h1e == _T_547 ? 8'h72 : _GEN_2853; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2855 = 8'h1f == _T_547 ? 8'hc0 : _GEN_2854; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2856 = 8'h20 == _T_547 ? 8'hb7 : _GEN_2855; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2857 = 8'h21 == _T_547 ? 8'hfd : _GEN_2856; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2858 = 8'h22 == _T_547 ? 8'h93 : _GEN_2857; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2859 = 8'h23 == _T_547 ? 8'h26 : _GEN_2858; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2860 = 8'h24 == _T_547 ? 8'h36 : _GEN_2859; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2861 = 8'h25 == _T_547 ? 8'h3f : _GEN_2860; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2862 = 8'h26 == _T_547 ? 8'hf7 : _GEN_2861; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2863 = 8'h27 == _T_547 ? 8'hcc : _GEN_2862; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2864 = 8'h28 == _T_547 ? 8'h34 : _GEN_2863; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2865 = 8'h29 == _T_547 ? 8'ha5 : _GEN_2864; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2866 = 8'h2a == _T_547 ? 8'he5 : _GEN_2865; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2867 = 8'h2b == _T_547 ? 8'hf1 : _GEN_2866; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2868 = 8'h2c == _T_547 ? 8'h71 : _GEN_2867; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2869 = 8'h2d == _T_547 ? 8'hd8 : _GEN_2868; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2870 = 8'h2e == _T_547 ? 8'h31 : _GEN_2869; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2871 = 8'h2f == _T_547 ? 8'h15 : _GEN_2870; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2872 = 8'h30 == _T_547 ? 8'h4 : _GEN_2871; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2873 = 8'h31 == _T_547 ? 8'hc7 : _GEN_2872; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2874 = 8'h32 == _T_547 ? 8'h23 : _GEN_2873; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2875 = 8'h33 == _T_547 ? 8'hc3 : _GEN_2874; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2876 = 8'h34 == _T_547 ? 8'h18 : _GEN_2875; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2877 = 8'h35 == _T_547 ? 8'h96 : _GEN_2876; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2878 = 8'h36 == _T_547 ? 8'h5 : _GEN_2877; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2879 = 8'h37 == _T_547 ? 8'h9a : _GEN_2878; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2880 = 8'h38 == _T_547 ? 8'h7 : _GEN_2879; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2881 = 8'h39 == _T_547 ? 8'h12 : _GEN_2880; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2882 = 8'h3a == _T_547 ? 8'h80 : _GEN_2881; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2883 = 8'h3b == _T_547 ? 8'he2 : _GEN_2882; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2884 = 8'h3c == _T_547 ? 8'heb : _GEN_2883; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2885 = 8'h3d == _T_547 ? 8'h27 : _GEN_2884; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2886 = 8'h3e == _T_547 ? 8'hb2 : _GEN_2885; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2887 = 8'h3f == _T_547 ? 8'h75 : _GEN_2886; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2888 = 8'h40 == _T_547 ? 8'h9 : _GEN_2887; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2889 = 8'h41 == _T_547 ? 8'h83 : _GEN_2888; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2890 = 8'h42 == _T_547 ? 8'h2c : _GEN_2889; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2891 = 8'h43 == _T_547 ? 8'h1a : _GEN_2890; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2892 = 8'h44 == _T_547 ? 8'h1b : _GEN_2891; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2893 = 8'h45 == _T_547 ? 8'h6e : _GEN_2892; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2894 = 8'h46 == _T_547 ? 8'h5a : _GEN_2893; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2895 = 8'h47 == _T_547 ? 8'ha0 : _GEN_2894; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2896 = 8'h48 == _T_547 ? 8'h52 : _GEN_2895; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2897 = 8'h49 == _T_547 ? 8'h3b : _GEN_2896; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2898 = 8'h4a == _T_547 ? 8'hd6 : _GEN_2897; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2899 = 8'h4b == _T_547 ? 8'hb3 : _GEN_2898; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2900 = 8'h4c == _T_547 ? 8'h29 : _GEN_2899; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2901 = 8'h4d == _T_547 ? 8'he3 : _GEN_2900; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2902 = 8'h4e == _T_547 ? 8'h2f : _GEN_2901; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2903 = 8'h4f == _T_547 ? 8'h84 : _GEN_2902; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2904 = 8'h50 == _T_547 ? 8'h53 : _GEN_2903; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2905 = 8'h51 == _T_547 ? 8'hd1 : _GEN_2904; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2906 = 8'h52 == _T_547 ? 8'h0 : _GEN_2905; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2907 = 8'h53 == _T_547 ? 8'hed : _GEN_2906; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2908 = 8'h54 == _T_547 ? 8'h20 : _GEN_2907; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2909 = 8'h55 == _T_547 ? 8'hfc : _GEN_2908; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2910 = 8'h56 == _T_547 ? 8'hb1 : _GEN_2909; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2911 = 8'h57 == _T_547 ? 8'h5b : _GEN_2910; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2912 = 8'h58 == _T_547 ? 8'h6a : _GEN_2911; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2913 = 8'h59 == _T_547 ? 8'hcb : _GEN_2912; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2914 = 8'h5a == _T_547 ? 8'hbe : _GEN_2913; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2915 = 8'h5b == _T_547 ? 8'h39 : _GEN_2914; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2916 = 8'h5c == _T_547 ? 8'h4a : _GEN_2915; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2917 = 8'h5d == _T_547 ? 8'h4c : _GEN_2916; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2918 = 8'h5e == _T_547 ? 8'h58 : _GEN_2917; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2919 = 8'h5f == _T_547 ? 8'hcf : _GEN_2918; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2920 = 8'h60 == _T_547 ? 8'hd0 : _GEN_2919; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2921 = 8'h61 == _T_547 ? 8'hef : _GEN_2920; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2922 = 8'h62 == _T_547 ? 8'haa : _GEN_2921; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2923 = 8'h63 == _T_547 ? 8'hfb : _GEN_2922; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2924 = 8'h64 == _T_547 ? 8'h43 : _GEN_2923; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2925 = 8'h65 == _T_547 ? 8'h4d : _GEN_2924; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2926 = 8'h66 == _T_547 ? 8'h33 : _GEN_2925; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2927 = 8'h67 == _T_547 ? 8'h85 : _GEN_2926; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2928 = 8'h68 == _T_547 ? 8'h45 : _GEN_2927; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2929 = 8'h69 == _T_547 ? 8'hf9 : _GEN_2928; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2930 = 8'h6a == _T_547 ? 8'h2 : _GEN_2929; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2931 = 8'h6b == _T_547 ? 8'h7f : _GEN_2930; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2932 = 8'h6c == _T_547 ? 8'h50 : _GEN_2931; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2933 = 8'h6d == _T_547 ? 8'h3c : _GEN_2932; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2934 = 8'h6e == _T_547 ? 8'h9f : _GEN_2933; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2935 = 8'h6f == _T_547 ? 8'ha8 : _GEN_2934; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2936 = 8'h70 == _T_547 ? 8'h51 : _GEN_2935; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2937 = 8'h71 == _T_547 ? 8'ha3 : _GEN_2936; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2938 = 8'h72 == _T_547 ? 8'h40 : _GEN_2937; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2939 = 8'h73 == _T_547 ? 8'h8f : _GEN_2938; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2940 = 8'h74 == _T_547 ? 8'h92 : _GEN_2939; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2941 = 8'h75 == _T_547 ? 8'h9d : _GEN_2940; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2942 = 8'h76 == _T_547 ? 8'h38 : _GEN_2941; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2943 = 8'h77 == _T_547 ? 8'hf5 : _GEN_2942; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2944 = 8'h78 == _T_547 ? 8'hbc : _GEN_2943; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2945 = 8'h79 == _T_547 ? 8'hb6 : _GEN_2944; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2946 = 8'h7a == _T_547 ? 8'hda : _GEN_2945; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2947 = 8'h7b == _T_547 ? 8'h21 : _GEN_2946; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2948 = 8'h7c == _T_547 ? 8'h10 : _GEN_2947; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2949 = 8'h7d == _T_547 ? 8'hff : _GEN_2948; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2950 = 8'h7e == _T_547 ? 8'hf3 : _GEN_2949; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2951 = 8'h7f == _T_547 ? 8'hd2 : _GEN_2950; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2952 = 8'h80 == _T_547 ? 8'hcd : _GEN_2951; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2953 = 8'h81 == _T_547 ? 8'hc : _GEN_2952; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2954 = 8'h82 == _T_547 ? 8'h13 : _GEN_2953; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2955 = 8'h83 == _T_547 ? 8'hec : _GEN_2954; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2956 = 8'h84 == _T_547 ? 8'h5f : _GEN_2955; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2957 = 8'h85 == _T_547 ? 8'h97 : _GEN_2956; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2958 = 8'h86 == _T_547 ? 8'h44 : _GEN_2957; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2959 = 8'h87 == _T_547 ? 8'h17 : _GEN_2958; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2960 = 8'h88 == _T_547 ? 8'hc4 : _GEN_2959; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2961 = 8'h89 == _T_547 ? 8'ha7 : _GEN_2960; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2962 = 8'h8a == _T_547 ? 8'h7e : _GEN_2961; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2963 = 8'h8b == _T_547 ? 8'h3d : _GEN_2962; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2964 = 8'h8c == _T_547 ? 8'h64 : _GEN_2963; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2965 = 8'h8d == _T_547 ? 8'h5d : _GEN_2964; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2966 = 8'h8e == _T_547 ? 8'h19 : _GEN_2965; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2967 = 8'h8f == _T_547 ? 8'h73 : _GEN_2966; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2968 = 8'h90 == _T_547 ? 8'h60 : _GEN_2967; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2969 = 8'h91 == _T_547 ? 8'h81 : _GEN_2968; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2970 = 8'h92 == _T_547 ? 8'h4f : _GEN_2969; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2971 = 8'h93 == _T_547 ? 8'hdc : _GEN_2970; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2972 = 8'h94 == _T_547 ? 8'h22 : _GEN_2971; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2973 = 8'h95 == _T_547 ? 8'h2a : _GEN_2972; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2974 = 8'h96 == _T_547 ? 8'h90 : _GEN_2973; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2975 = 8'h97 == _T_547 ? 8'h88 : _GEN_2974; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2976 = 8'h98 == _T_547 ? 8'h46 : _GEN_2975; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2977 = 8'h99 == _T_547 ? 8'hee : _GEN_2976; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2978 = 8'h9a == _T_547 ? 8'hb8 : _GEN_2977; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2979 = 8'h9b == _T_547 ? 8'h14 : _GEN_2978; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2980 = 8'h9c == _T_547 ? 8'hde : _GEN_2979; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2981 = 8'h9d == _T_547 ? 8'h5e : _GEN_2980; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2982 = 8'h9e == _T_547 ? 8'hb : _GEN_2981; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2983 = 8'h9f == _T_547 ? 8'hdb : _GEN_2982; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2984 = 8'ha0 == _T_547 ? 8'he0 : _GEN_2983; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2985 = 8'ha1 == _T_547 ? 8'h32 : _GEN_2984; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2986 = 8'ha2 == _T_547 ? 8'h3a : _GEN_2985; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2987 = 8'ha3 == _T_547 ? 8'ha : _GEN_2986; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2988 = 8'ha4 == _T_547 ? 8'h49 : _GEN_2987; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2989 = 8'ha5 == _T_547 ? 8'h6 : _GEN_2988; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2990 = 8'ha6 == _T_547 ? 8'h24 : _GEN_2989; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2991 = 8'ha7 == _T_547 ? 8'h5c : _GEN_2990; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2992 = 8'ha8 == _T_547 ? 8'hc2 : _GEN_2991; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2993 = 8'ha9 == _T_547 ? 8'hd3 : _GEN_2992; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2994 = 8'haa == _T_547 ? 8'hac : _GEN_2993; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2995 = 8'hab == _T_547 ? 8'h62 : _GEN_2994; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2996 = 8'hac == _T_547 ? 8'h91 : _GEN_2995; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2997 = 8'had == _T_547 ? 8'h95 : _GEN_2996; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2998 = 8'hae == _T_547 ? 8'he4 : _GEN_2997; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_2999 = 8'haf == _T_547 ? 8'h79 : _GEN_2998; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3000 = 8'hb0 == _T_547 ? 8'he7 : _GEN_2999; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3001 = 8'hb1 == _T_547 ? 8'hc8 : _GEN_3000; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3002 = 8'hb2 == _T_547 ? 8'h37 : _GEN_3001; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3003 = 8'hb3 == _T_547 ? 8'h6d : _GEN_3002; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3004 = 8'hb4 == _T_547 ? 8'h8d : _GEN_3003; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3005 = 8'hb5 == _T_547 ? 8'hd5 : _GEN_3004; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3006 = 8'hb6 == _T_547 ? 8'h4e : _GEN_3005; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3007 = 8'hb7 == _T_547 ? 8'ha9 : _GEN_3006; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3008 = 8'hb8 == _T_547 ? 8'h6c : _GEN_3007; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3009 = 8'hb9 == _T_547 ? 8'h56 : _GEN_3008; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3010 = 8'hba == _T_547 ? 8'hf4 : _GEN_3009; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3011 = 8'hbb == _T_547 ? 8'hea : _GEN_3010; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3012 = 8'hbc == _T_547 ? 8'h65 : _GEN_3011; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3013 = 8'hbd == _T_547 ? 8'h7a : _GEN_3012; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3014 = 8'hbe == _T_547 ? 8'hae : _GEN_3013; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3015 = 8'hbf == _T_547 ? 8'h8 : _GEN_3014; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3016 = 8'hc0 == _T_547 ? 8'hba : _GEN_3015; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3017 = 8'hc1 == _T_547 ? 8'h78 : _GEN_3016; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3018 = 8'hc2 == _T_547 ? 8'h25 : _GEN_3017; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3019 = 8'hc3 == _T_547 ? 8'h2e : _GEN_3018; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3020 = 8'hc4 == _T_547 ? 8'h1c : _GEN_3019; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3021 = 8'hc5 == _T_547 ? 8'ha6 : _GEN_3020; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3022 = 8'hc6 == _T_547 ? 8'hb4 : _GEN_3021; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3023 = 8'hc7 == _T_547 ? 8'hc6 : _GEN_3022; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3024 = 8'hc8 == _T_547 ? 8'he8 : _GEN_3023; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3025 = 8'hc9 == _T_547 ? 8'hdd : _GEN_3024; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3026 = 8'hca == _T_547 ? 8'h74 : _GEN_3025; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3027 = 8'hcb == _T_547 ? 8'h1f : _GEN_3026; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3028 = 8'hcc == _T_547 ? 8'h4b : _GEN_3027; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3029 = 8'hcd == _T_547 ? 8'hbd : _GEN_3028; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3030 = 8'hce == _T_547 ? 8'h8b : _GEN_3029; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3031 = 8'hcf == _T_547 ? 8'h8a : _GEN_3030; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3032 = 8'hd0 == _T_547 ? 8'h70 : _GEN_3031; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3033 = 8'hd1 == _T_547 ? 8'h3e : _GEN_3032; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3034 = 8'hd2 == _T_547 ? 8'hb5 : _GEN_3033; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3035 = 8'hd3 == _T_547 ? 8'h66 : _GEN_3034; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3036 = 8'hd4 == _T_547 ? 8'h48 : _GEN_3035; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3037 = 8'hd5 == _T_547 ? 8'h3 : _GEN_3036; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3038 = 8'hd6 == _T_547 ? 8'hf6 : _GEN_3037; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3039 = 8'hd7 == _T_547 ? 8'he : _GEN_3038; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3040 = 8'hd8 == _T_547 ? 8'h61 : _GEN_3039; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3041 = 8'hd9 == _T_547 ? 8'h35 : _GEN_3040; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3042 = 8'hda == _T_547 ? 8'h57 : _GEN_3041; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3043 = 8'hdb == _T_547 ? 8'hb9 : _GEN_3042; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3044 = 8'hdc == _T_547 ? 8'h86 : _GEN_3043; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3045 = 8'hdd == _T_547 ? 8'hc1 : _GEN_3044; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3046 = 8'hde == _T_547 ? 8'h1d : _GEN_3045; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3047 = 8'hdf == _T_547 ? 8'h9e : _GEN_3046; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3048 = 8'he0 == _T_547 ? 8'he1 : _GEN_3047; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3049 = 8'he1 == _T_547 ? 8'hf8 : _GEN_3048; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3050 = 8'he2 == _T_547 ? 8'h98 : _GEN_3049; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3051 = 8'he3 == _T_547 ? 8'h11 : _GEN_3050; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3052 = 8'he4 == _T_547 ? 8'h69 : _GEN_3051; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3053 = 8'he5 == _T_547 ? 8'hd9 : _GEN_3052; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3054 = 8'he6 == _T_547 ? 8'h8e : _GEN_3053; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3055 = 8'he7 == _T_547 ? 8'h94 : _GEN_3054; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3056 = 8'he8 == _T_547 ? 8'h9b : _GEN_3055; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3057 = 8'he9 == _T_547 ? 8'h1e : _GEN_3056; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3058 = 8'hea == _T_547 ? 8'h87 : _GEN_3057; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3059 = 8'heb == _T_547 ? 8'he9 : _GEN_3058; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3060 = 8'hec == _T_547 ? 8'hce : _GEN_3059; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3061 = 8'hed == _T_547 ? 8'h55 : _GEN_3060; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3062 = 8'hee == _T_547 ? 8'h28 : _GEN_3061; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3063 = 8'hef == _T_547 ? 8'hdf : _GEN_3062; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3064 = 8'hf0 == _T_547 ? 8'h8c : _GEN_3063; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3065 = 8'hf1 == _T_547 ? 8'ha1 : _GEN_3064; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3066 = 8'hf2 == _T_547 ? 8'h89 : _GEN_3065; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3067 = 8'hf3 == _T_547 ? 8'hd : _GEN_3066; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3068 = 8'hf4 == _T_547 ? 8'hbf : _GEN_3067; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3069 = 8'hf5 == _T_547 ? 8'he6 : _GEN_3068; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3070 = 8'hf6 == _T_547 ? 8'h42 : _GEN_3069; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3071 = 8'hf7 == _T_547 ? 8'h68 : _GEN_3070; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3072 = 8'hf8 == _T_547 ? 8'h41 : _GEN_3071; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3073 = 8'hf9 == _T_547 ? 8'h99 : _GEN_3072; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3074 = 8'hfa == _T_547 ? 8'h2d : _GEN_3073; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3075 = 8'hfb == _T_547 ? 8'hf : _GEN_3074; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3076 = 8'hfc == _T_547 ? 8'hb0 : _GEN_3075; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3077 = 8'hfd == _T_547 ? 8'h54 : _GEN_3076; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3078 = 8'hfe == _T_547 ? 8'hbb : _GEN_3077; // @[Cat.scala 30:58:@2081.4]
  assign _GEN_3079 = 8'hff == _T_547 ? 8'h16 : _GEN_3078; // @[Cat.scala 30:58:@2081.4]
  assign _T_552 = {_GEN_2824,_GEN_3079}; // @[Cat.scala 30:58:@2081.4]
  assign x2 = {_T_552,_T_551}; // @[Cat.scala 30:58:@2082.4]
  assign _T_553 = io_addr2[71:64]; // @[sbox.scala 69:26:@2083.4]
  assign _T_555 = io_addr2[79:72]; // @[sbox.scala 70:26:@2084.4]
  assign _T_557 = io_addr2[87:80]; // @[sbox.scala 71:26:@2085.4]
  assign _T_559 = io_addr2[95:88]; // @[sbox.scala 72:26:@2086.4]
  assign _GEN_3080 = 8'h1 == _T_555 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3081 = 8'h2 == _T_555 ? 8'h77 : _GEN_3080; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3082 = 8'h3 == _T_555 ? 8'h7b : _GEN_3081; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3083 = 8'h4 == _T_555 ? 8'hf2 : _GEN_3082; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3084 = 8'h5 == _T_555 ? 8'h6b : _GEN_3083; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3085 = 8'h6 == _T_555 ? 8'h6f : _GEN_3084; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3086 = 8'h7 == _T_555 ? 8'hc5 : _GEN_3085; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3087 = 8'h8 == _T_555 ? 8'h30 : _GEN_3086; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3088 = 8'h9 == _T_555 ? 8'h1 : _GEN_3087; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3089 = 8'ha == _T_555 ? 8'h67 : _GEN_3088; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3090 = 8'hb == _T_555 ? 8'h2b : _GEN_3089; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3091 = 8'hc == _T_555 ? 8'hfe : _GEN_3090; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3092 = 8'hd == _T_555 ? 8'hd7 : _GEN_3091; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3093 = 8'he == _T_555 ? 8'hab : _GEN_3092; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3094 = 8'hf == _T_555 ? 8'h76 : _GEN_3093; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3095 = 8'h10 == _T_555 ? 8'hca : _GEN_3094; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3096 = 8'h11 == _T_555 ? 8'h82 : _GEN_3095; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3097 = 8'h12 == _T_555 ? 8'hc9 : _GEN_3096; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3098 = 8'h13 == _T_555 ? 8'h7d : _GEN_3097; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3099 = 8'h14 == _T_555 ? 8'hfa : _GEN_3098; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3100 = 8'h15 == _T_555 ? 8'h59 : _GEN_3099; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3101 = 8'h16 == _T_555 ? 8'h47 : _GEN_3100; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3102 = 8'h17 == _T_555 ? 8'hf0 : _GEN_3101; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3103 = 8'h18 == _T_555 ? 8'had : _GEN_3102; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3104 = 8'h19 == _T_555 ? 8'hd4 : _GEN_3103; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3105 = 8'h1a == _T_555 ? 8'ha2 : _GEN_3104; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3106 = 8'h1b == _T_555 ? 8'haf : _GEN_3105; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3107 = 8'h1c == _T_555 ? 8'h9c : _GEN_3106; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3108 = 8'h1d == _T_555 ? 8'ha4 : _GEN_3107; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3109 = 8'h1e == _T_555 ? 8'h72 : _GEN_3108; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3110 = 8'h1f == _T_555 ? 8'hc0 : _GEN_3109; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3111 = 8'h20 == _T_555 ? 8'hb7 : _GEN_3110; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3112 = 8'h21 == _T_555 ? 8'hfd : _GEN_3111; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3113 = 8'h22 == _T_555 ? 8'h93 : _GEN_3112; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3114 = 8'h23 == _T_555 ? 8'h26 : _GEN_3113; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3115 = 8'h24 == _T_555 ? 8'h36 : _GEN_3114; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3116 = 8'h25 == _T_555 ? 8'h3f : _GEN_3115; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3117 = 8'h26 == _T_555 ? 8'hf7 : _GEN_3116; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3118 = 8'h27 == _T_555 ? 8'hcc : _GEN_3117; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3119 = 8'h28 == _T_555 ? 8'h34 : _GEN_3118; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3120 = 8'h29 == _T_555 ? 8'ha5 : _GEN_3119; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3121 = 8'h2a == _T_555 ? 8'he5 : _GEN_3120; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3122 = 8'h2b == _T_555 ? 8'hf1 : _GEN_3121; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3123 = 8'h2c == _T_555 ? 8'h71 : _GEN_3122; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3124 = 8'h2d == _T_555 ? 8'hd8 : _GEN_3123; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3125 = 8'h2e == _T_555 ? 8'h31 : _GEN_3124; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3126 = 8'h2f == _T_555 ? 8'h15 : _GEN_3125; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3127 = 8'h30 == _T_555 ? 8'h4 : _GEN_3126; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3128 = 8'h31 == _T_555 ? 8'hc7 : _GEN_3127; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3129 = 8'h32 == _T_555 ? 8'h23 : _GEN_3128; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3130 = 8'h33 == _T_555 ? 8'hc3 : _GEN_3129; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3131 = 8'h34 == _T_555 ? 8'h18 : _GEN_3130; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3132 = 8'h35 == _T_555 ? 8'h96 : _GEN_3131; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3133 = 8'h36 == _T_555 ? 8'h5 : _GEN_3132; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3134 = 8'h37 == _T_555 ? 8'h9a : _GEN_3133; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3135 = 8'h38 == _T_555 ? 8'h7 : _GEN_3134; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3136 = 8'h39 == _T_555 ? 8'h12 : _GEN_3135; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3137 = 8'h3a == _T_555 ? 8'h80 : _GEN_3136; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3138 = 8'h3b == _T_555 ? 8'he2 : _GEN_3137; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3139 = 8'h3c == _T_555 ? 8'heb : _GEN_3138; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3140 = 8'h3d == _T_555 ? 8'h27 : _GEN_3139; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3141 = 8'h3e == _T_555 ? 8'hb2 : _GEN_3140; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3142 = 8'h3f == _T_555 ? 8'h75 : _GEN_3141; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3143 = 8'h40 == _T_555 ? 8'h9 : _GEN_3142; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3144 = 8'h41 == _T_555 ? 8'h83 : _GEN_3143; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3145 = 8'h42 == _T_555 ? 8'h2c : _GEN_3144; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3146 = 8'h43 == _T_555 ? 8'h1a : _GEN_3145; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3147 = 8'h44 == _T_555 ? 8'h1b : _GEN_3146; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3148 = 8'h45 == _T_555 ? 8'h6e : _GEN_3147; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3149 = 8'h46 == _T_555 ? 8'h5a : _GEN_3148; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3150 = 8'h47 == _T_555 ? 8'ha0 : _GEN_3149; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3151 = 8'h48 == _T_555 ? 8'h52 : _GEN_3150; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3152 = 8'h49 == _T_555 ? 8'h3b : _GEN_3151; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3153 = 8'h4a == _T_555 ? 8'hd6 : _GEN_3152; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3154 = 8'h4b == _T_555 ? 8'hb3 : _GEN_3153; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3155 = 8'h4c == _T_555 ? 8'h29 : _GEN_3154; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3156 = 8'h4d == _T_555 ? 8'he3 : _GEN_3155; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3157 = 8'h4e == _T_555 ? 8'h2f : _GEN_3156; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3158 = 8'h4f == _T_555 ? 8'h84 : _GEN_3157; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3159 = 8'h50 == _T_555 ? 8'h53 : _GEN_3158; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3160 = 8'h51 == _T_555 ? 8'hd1 : _GEN_3159; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3161 = 8'h52 == _T_555 ? 8'h0 : _GEN_3160; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3162 = 8'h53 == _T_555 ? 8'hed : _GEN_3161; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3163 = 8'h54 == _T_555 ? 8'h20 : _GEN_3162; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3164 = 8'h55 == _T_555 ? 8'hfc : _GEN_3163; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3165 = 8'h56 == _T_555 ? 8'hb1 : _GEN_3164; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3166 = 8'h57 == _T_555 ? 8'h5b : _GEN_3165; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3167 = 8'h58 == _T_555 ? 8'h6a : _GEN_3166; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3168 = 8'h59 == _T_555 ? 8'hcb : _GEN_3167; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3169 = 8'h5a == _T_555 ? 8'hbe : _GEN_3168; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3170 = 8'h5b == _T_555 ? 8'h39 : _GEN_3169; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3171 = 8'h5c == _T_555 ? 8'h4a : _GEN_3170; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3172 = 8'h5d == _T_555 ? 8'h4c : _GEN_3171; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3173 = 8'h5e == _T_555 ? 8'h58 : _GEN_3172; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3174 = 8'h5f == _T_555 ? 8'hcf : _GEN_3173; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3175 = 8'h60 == _T_555 ? 8'hd0 : _GEN_3174; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3176 = 8'h61 == _T_555 ? 8'hef : _GEN_3175; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3177 = 8'h62 == _T_555 ? 8'haa : _GEN_3176; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3178 = 8'h63 == _T_555 ? 8'hfb : _GEN_3177; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3179 = 8'h64 == _T_555 ? 8'h43 : _GEN_3178; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3180 = 8'h65 == _T_555 ? 8'h4d : _GEN_3179; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3181 = 8'h66 == _T_555 ? 8'h33 : _GEN_3180; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3182 = 8'h67 == _T_555 ? 8'h85 : _GEN_3181; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3183 = 8'h68 == _T_555 ? 8'h45 : _GEN_3182; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3184 = 8'h69 == _T_555 ? 8'hf9 : _GEN_3183; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3185 = 8'h6a == _T_555 ? 8'h2 : _GEN_3184; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3186 = 8'h6b == _T_555 ? 8'h7f : _GEN_3185; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3187 = 8'h6c == _T_555 ? 8'h50 : _GEN_3186; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3188 = 8'h6d == _T_555 ? 8'h3c : _GEN_3187; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3189 = 8'h6e == _T_555 ? 8'h9f : _GEN_3188; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3190 = 8'h6f == _T_555 ? 8'ha8 : _GEN_3189; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3191 = 8'h70 == _T_555 ? 8'h51 : _GEN_3190; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3192 = 8'h71 == _T_555 ? 8'ha3 : _GEN_3191; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3193 = 8'h72 == _T_555 ? 8'h40 : _GEN_3192; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3194 = 8'h73 == _T_555 ? 8'h8f : _GEN_3193; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3195 = 8'h74 == _T_555 ? 8'h92 : _GEN_3194; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3196 = 8'h75 == _T_555 ? 8'h9d : _GEN_3195; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3197 = 8'h76 == _T_555 ? 8'h38 : _GEN_3196; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3198 = 8'h77 == _T_555 ? 8'hf5 : _GEN_3197; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3199 = 8'h78 == _T_555 ? 8'hbc : _GEN_3198; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3200 = 8'h79 == _T_555 ? 8'hb6 : _GEN_3199; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3201 = 8'h7a == _T_555 ? 8'hda : _GEN_3200; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3202 = 8'h7b == _T_555 ? 8'h21 : _GEN_3201; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3203 = 8'h7c == _T_555 ? 8'h10 : _GEN_3202; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3204 = 8'h7d == _T_555 ? 8'hff : _GEN_3203; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3205 = 8'h7e == _T_555 ? 8'hf3 : _GEN_3204; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3206 = 8'h7f == _T_555 ? 8'hd2 : _GEN_3205; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3207 = 8'h80 == _T_555 ? 8'hcd : _GEN_3206; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3208 = 8'h81 == _T_555 ? 8'hc : _GEN_3207; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3209 = 8'h82 == _T_555 ? 8'h13 : _GEN_3208; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3210 = 8'h83 == _T_555 ? 8'hec : _GEN_3209; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3211 = 8'h84 == _T_555 ? 8'h5f : _GEN_3210; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3212 = 8'h85 == _T_555 ? 8'h97 : _GEN_3211; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3213 = 8'h86 == _T_555 ? 8'h44 : _GEN_3212; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3214 = 8'h87 == _T_555 ? 8'h17 : _GEN_3213; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3215 = 8'h88 == _T_555 ? 8'hc4 : _GEN_3214; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3216 = 8'h89 == _T_555 ? 8'ha7 : _GEN_3215; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3217 = 8'h8a == _T_555 ? 8'h7e : _GEN_3216; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3218 = 8'h8b == _T_555 ? 8'h3d : _GEN_3217; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3219 = 8'h8c == _T_555 ? 8'h64 : _GEN_3218; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3220 = 8'h8d == _T_555 ? 8'h5d : _GEN_3219; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3221 = 8'h8e == _T_555 ? 8'h19 : _GEN_3220; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3222 = 8'h8f == _T_555 ? 8'h73 : _GEN_3221; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3223 = 8'h90 == _T_555 ? 8'h60 : _GEN_3222; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3224 = 8'h91 == _T_555 ? 8'h81 : _GEN_3223; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3225 = 8'h92 == _T_555 ? 8'h4f : _GEN_3224; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3226 = 8'h93 == _T_555 ? 8'hdc : _GEN_3225; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3227 = 8'h94 == _T_555 ? 8'h22 : _GEN_3226; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3228 = 8'h95 == _T_555 ? 8'h2a : _GEN_3227; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3229 = 8'h96 == _T_555 ? 8'h90 : _GEN_3228; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3230 = 8'h97 == _T_555 ? 8'h88 : _GEN_3229; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3231 = 8'h98 == _T_555 ? 8'h46 : _GEN_3230; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3232 = 8'h99 == _T_555 ? 8'hee : _GEN_3231; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3233 = 8'h9a == _T_555 ? 8'hb8 : _GEN_3232; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3234 = 8'h9b == _T_555 ? 8'h14 : _GEN_3233; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3235 = 8'h9c == _T_555 ? 8'hde : _GEN_3234; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3236 = 8'h9d == _T_555 ? 8'h5e : _GEN_3235; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3237 = 8'h9e == _T_555 ? 8'hb : _GEN_3236; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3238 = 8'h9f == _T_555 ? 8'hdb : _GEN_3237; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3239 = 8'ha0 == _T_555 ? 8'he0 : _GEN_3238; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3240 = 8'ha1 == _T_555 ? 8'h32 : _GEN_3239; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3241 = 8'ha2 == _T_555 ? 8'h3a : _GEN_3240; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3242 = 8'ha3 == _T_555 ? 8'ha : _GEN_3241; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3243 = 8'ha4 == _T_555 ? 8'h49 : _GEN_3242; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3244 = 8'ha5 == _T_555 ? 8'h6 : _GEN_3243; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3245 = 8'ha6 == _T_555 ? 8'h24 : _GEN_3244; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3246 = 8'ha7 == _T_555 ? 8'h5c : _GEN_3245; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3247 = 8'ha8 == _T_555 ? 8'hc2 : _GEN_3246; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3248 = 8'ha9 == _T_555 ? 8'hd3 : _GEN_3247; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3249 = 8'haa == _T_555 ? 8'hac : _GEN_3248; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3250 = 8'hab == _T_555 ? 8'h62 : _GEN_3249; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3251 = 8'hac == _T_555 ? 8'h91 : _GEN_3250; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3252 = 8'had == _T_555 ? 8'h95 : _GEN_3251; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3253 = 8'hae == _T_555 ? 8'he4 : _GEN_3252; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3254 = 8'haf == _T_555 ? 8'h79 : _GEN_3253; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3255 = 8'hb0 == _T_555 ? 8'he7 : _GEN_3254; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3256 = 8'hb1 == _T_555 ? 8'hc8 : _GEN_3255; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3257 = 8'hb2 == _T_555 ? 8'h37 : _GEN_3256; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3258 = 8'hb3 == _T_555 ? 8'h6d : _GEN_3257; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3259 = 8'hb4 == _T_555 ? 8'h8d : _GEN_3258; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3260 = 8'hb5 == _T_555 ? 8'hd5 : _GEN_3259; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3261 = 8'hb6 == _T_555 ? 8'h4e : _GEN_3260; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3262 = 8'hb7 == _T_555 ? 8'ha9 : _GEN_3261; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3263 = 8'hb8 == _T_555 ? 8'h6c : _GEN_3262; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3264 = 8'hb9 == _T_555 ? 8'h56 : _GEN_3263; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3265 = 8'hba == _T_555 ? 8'hf4 : _GEN_3264; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3266 = 8'hbb == _T_555 ? 8'hea : _GEN_3265; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3267 = 8'hbc == _T_555 ? 8'h65 : _GEN_3266; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3268 = 8'hbd == _T_555 ? 8'h7a : _GEN_3267; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3269 = 8'hbe == _T_555 ? 8'hae : _GEN_3268; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3270 = 8'hbf == _T_555 ? 8'h8 : _GEN_3269; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3271 = 8'hc0 == _T_555 ? 8'hba : _GEN_3270; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3272 = 8'hc1 == _T_555 ? 8'h78 : _GEN_3271; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3273 = 8'hc2 == _T_555 ? 8'h25 : _GEN_3272; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3274 = 8'hc3 == _T_555 ? 8'h2e : _GEN_3273; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3275 = 8'hc4 == _T_555 ? 8'h1c : _GEN_3274; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3276 = 8'hc5 == _T_555 ? 8'ha6 : _GEN_3275; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3277 = 8'hc6 == _T_555 ? 8'hb4 : _GEN_3276; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3278 = 8'hc7 == _T_555 ? 8'hc6 : _GEN_3277; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3279 = 8'hc8 == _T_555 ? 8'he8 : _GEN_3278; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3280 = 8'hc9 == _T_555 ? 8'hdd : _GEN_3279; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3281 = 8'hca == _T_555 ? 8'h74 : _GEN_3280; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3282 = 8'hcb == _T_555 ? 8'h1f : _GEN_3281; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3283 = 8'hcc == _T_555 ? 8'h4b : _GEN_3282; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3284 = 8'hcd == _T_555 ? 8'hbd : _GEN_3283; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3285 = 8'hce == _T_555 ? 8'h8b : _GEN_3284; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3286 = 8'hcf == _T_555 ? 8'h8a : _GEN_3285; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3287 = 8'hd0 == _T_555 ? 8'h70 : _GEN_3286; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3288 = 8'hd1 == _T_555 ? 8'h3e : _GEN_3287; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3289 = 8'hd2 == _T_555 ? 8'hb5 : _GEN_3288; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3290 = 8'hd3 == _T_555 ? 8'h66 : _GEN_3289; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3291 = 8'hd4 == _T_555 ? 8'h48 : _GEN_3290; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3292 = 8'hd5 == _T_555 ? 8'h3 : _GEN_3291; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3293 = 8'hd6 == _T_555 ? 8'hf6 : _GEN_3292; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3294 = 8'hd7 == _T_555 ? 8'he : _GEN_3293; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3295 = 8'hd8 == _T_555 ? 8'h61 : _GEN_3294; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3296 = 8'hd9 == _T_555 ? 8'h35 : _GEN_3295; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3297 = 8'hda == _T_555 ? 8'h57 : _GEN_3296; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3298 = 8'hdb == _T_555 ? 8'hb9 : _GEN_3297; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3299 = 8'hdc == _T_555 ? 8'h86 : _GEN_3298; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3300 = 8'hdd == _T_555 ? 8'hc1 : _GEN_3299; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3301 = 8'hde == _T_555 ? 8'h1d : _GEN_3300; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3302 = 8'hdf == _T_555 ? 8'h9e : _GEN_3301; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3303 = 8'he0 == _T_555 ? 8'he1 : _GEN_3302; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3304 = 8'he1 == _T_555 ? 8'hf8 : _GEN_3303; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3305 = 8'he2 == _T_555 ? 8'h98 : _GEN_3304; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3306 = 8'he3 == _T_555 ? 8'h11 : _GEN_3305; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3307 = 8'he4 == _T_555 ? 8'h69 : _GEN_3306; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3308 = 8'he5 == _T_555 ? 8'hd9 : _GEN_3307; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3309 = 8'he6 == _T_555 ? 8'h8e : _GEN_3308; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3310 = 8'he7 == _T_555 ? 8'h94 : _GEN_3309; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3311 = 8'he8 == _T_555 ? 8'h9b : _GEN_3310; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3312 = 8'he9 == _T_555 ? 8'h1e : _GEN_3311; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3313 = 8'hea == _T_555 ? 8'h87 : _GEN_3312; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3314 = 8'heb == _T_555 ? 8'he9 : _GEN_3313; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3315 = 8'hec == _T_555 ? 8'hce : _GEN_3314; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3316 = 8'hed == _T_555 ? 8'h55 : _GEN_3315; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3317 = 8'hee == _T_555 ? 8'h28 : _GEN_3316; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3318 = 8'hef == _T_555 ? 8'hdf : _GEN_3317; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3319 = 8'hf0 == _T_555 ? 8'h8c : _GEN_3318; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3320 = 8'hf1 == _T_555 ? 8'ha1 : _GEN_3319; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3321 = 8'hf2 == _T_555 ? 8'h89 : _GEN_3320; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3322 = 8'hf3 == _T_555 ? 8'hd : _GEN_3321; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3323 = 8'hf4 == _T_555 ? 8'hbf : _GEN_3322; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3324 = 8'hf5 == _T_555 ? 8'he6 : _GEN_3323; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3325 = 8'hf6 == _T_555 ? 8'h42 : _GEN_3324; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3326 = 8'hf7 == _T_555 ? 8'h68 : _GEN_3325; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3327 = 8'hf8 == _T_555 ? 8'h41 : _GEN_3326; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3328 = 8'hf9 == _T_555 ? 8'h99 : _GEN_3327; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3329 = 8'hfa == _T_555 ? 8'h2d : _GEN_3328; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3330 = 8'hfb == _T_555 ? 8'hf : _GEN_3329; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3331 = 8'hfc == _T_555 ? 8'hb0 : _GEN_3330; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3332 = 8'hfd == _T_555 ? 8'h54 : _GEN_3331; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3333 = 8'hfe == _T_555 ? 8'hbb : _GEN_3332; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3334 = 8'hff == _T_555 ? 8'h16 : _GEN_3333; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3335 = 8'h1 == _T_553 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3336 = 8'h2 == _T_553 ? 8'h77 : _GEN_3335; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3337 = 8'h3 == _T_553 ? 8'h7b : _GEN_3336; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3338 = 8'h4 == _T_553 ? 8'hf2 : _GEN_3337; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3339 = 8'h5 == _T_553 ? 8'h6b : _GEN_3338; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3340 = 8'h6 == _T_553 ? 8'h6f : _GEN_3339; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3341 = 8'h7 == _T_553 ? 8'hc5 : _GEN_3340; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3342 = 8'h8 == _T_553 ? 8'h30 : _GEN_3341; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3343 = 8'h9 == _T_553 ? 8'h1 : _GEN_3342; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3344 = 8'ha == _T_553 ? 8'h67 : _GEN_3343; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3345 = 8'hb == _T_553 ? 8'h2b : _GEN_3344; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3346 = 8'hc == _T_553 ? 8'hfe : _GEN_3345; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3347 = 8'hd == _T_553 ? 8'hd7 : _GEN_3346; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3348 = 8'he == _T_553 ? 8'hab : _GEN_3347; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3349 = 8'hf == _T_553 ? 8'h76 : _GEN_3348; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3350 = 8'h10 == _T_553 ? 8'hca : _GEN_3349; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3351 = 8'h11 == _T_553 ? 8'h82 : _GEN_3350; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3352 = 8'h12 == _T_553 ? 8'hc9 : _GEN_3351; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3353 = 8'h13 == _T_553 ? 8'h7d : _GEN_3352; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3354 = 8'h14 == _T_553 ? 8'hfa : _GEN_3353; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3355 = 8'h15 == _T_553 ? 8'h59 : _GEN_3354; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3356 = 8'h16 == _T_553 ? 8'h47 : _GEN_3355; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3357 = 8'h17 == _T_553 ? 8'hf0 : _GEN_3356; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3358 = 8'h18 == _T_553 ? 8'had : _GEN_3357; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3359 = 8'h19 == _T_553 ? 8'hd4 : _GEN_3358; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3360 = 8'h1a == _T_553 ? 8'ha2 : _GEN_3359; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3361 = 8'h1b == _T_553 ? 8'haf : _GEN_3360; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3362 = 8'h1c == _T_553 ? 8'h9c : _GEN_3361; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3363 = 8'h1d == _T_553 ? 8'ha4 : _GEN_3362; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3364 = 8'h1e == _T_553 ? 8'h72 : _GEN_3363; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3365 = 8'h1f == _T_553 ? 8'hc0 : _GEN_3364; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3366 = 8'h20 == _T_553 ? 8'hb7 : _GEN_3365; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3367 = 8'h21 == _T_553 ? 8'hfd : _GEN_3366; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3368 = 8'h22 == _T_553 ? 8'h93 : _GEN_3367; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3369 = 8'h23 == _T_553 ? 8'h26 : _GEN_3368; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3370 = 8'h24 == _T_553 ? 8'h36 : _GEN_3369; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3371 = 8'h25 == _T_553 ? 8'h3f : _GEN_3370; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3372 = 8'h26 == _T_553 ? 8'hf7 : _GEN_3371; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3373 = 8'h27 == _T_553 ? 8'hcc : _GEN_3372; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3374 = 8'h28 == _T_553 ? 8'h34 : _GEN_3373; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3375 = 8'h29 == _T_553 ? 8'ha5 : _GEN_3374; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3376 = 8'h2a == _T_553 ? 8'he5 : _GEN_3375; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3377 = 8'h2b == _T_553 ? 8'hf1 : _GEN_3376; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3378 = 8'h2c == _T_553 ? 8'h71 : _GEN_3377; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3379 = 8'h2d == _T_553 ? 8'hd8 : _GEN_3378; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3380 = 8'h2e == _T_553 ? 8'h31 : _GEN_3379; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3381 = 8'h2f == _T_553 ? 8'h15 : _GEN_3380; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3382 = 8'h30 == _T_553 ? 8'h4 : _GEN_3381; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3383 = 8'h31 == _T_553 ? 8'hc7 : _GEN_3382; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3384 = 8'h32 == _T_553 ? 8'h23 : _GEN_3383; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3385 = 8'h33 == _T_553 ? 8'hc3 : _GEN_3384; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3386 = 8'h34 == _T_553 ? 8'h18 : _GEN_3385; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3387 = 8'h35 == _T_553 ? 8'h96 : _GEN_3386; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3388 = 8'h36 == _T_553 ? 8'h5 : _GEN_3387; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3389 = 8'h37 == _T_553 ? 8'h9a : _GEN_3388; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3390 = 8'h38 == _T_553 ? 8'h7 : _GEN_3389; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3391 = 8'h39 == _T_553 ? 8'h12 : _GEN_3390; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3392 = 8'h3a == _T_553 ? 8'h80 : _GEN_3391; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3393 = 8'h3b == _T_553 ? 8'he2 : _GEN_3392; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3394 = 8'h3c == _T_553 ? 8'heb : _GEN_3393; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3395 = 8'h3d == _T_553 ? 8'h27 : _GEN_3394; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3396 = 8'h3e == _T_553 ? 8'hb2 : _GEN_3395; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3397 = 8'h3f == _T_553 ? 8'h75 : _GEN_3396; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3398 = 8'h40 == _T_553 ? 8'h9 : _GEN_3397; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3399 = 8'h41 == _T_553 ? 8'h83 : _GEN_3398; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3400 = 8'h42 == _T_553 ? 8'h2c : _GEN_3399; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3401 = 8'h43 == _T_553 ? 8'h1a : _GEN_3400; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3402 = 8'h44 == _T_553 ? 8'h1b : _GEN_3401; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3403 = 8'h45 == _T_553 ? 8'h6e : _GEN_3402; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3404 = 8'h46 == _T_553 ? 8'h5a : _GEN_3403; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3405 = 8'h47 == _T_553 ? 8'ha0 : _GEN_3404; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3406 = 8'h48 == _T_553 ? 8'h52 : _GEN_3405; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3407 = 8'h49 == _T_553 ? 8'h3b : _GEN_3406; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3408 = 8'h4a == _T_553 ? 8'hd6 : _GEN_3407; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3409 = 8'h4b == _T_553 ? 8'hb3 : _GEN_3408; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3410 = 8'h4c == _T_553 ? 8'h29 : _GEN_3409; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3411 = 8'h4d == _T_553 ? 8'he3 : _GEN_3410; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3412 = 8'h4e == _T_553 ? 8'h2f : _GEN_3411; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3413 = 8'h4f == _T_553 ? 8'h84 : _GEN_3412; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3414 = 8'h50 == _T_553 ? 8'h53 : _GEN_3413; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3415 = 8'h51 == _T_553 ? 8'hd1 : _GEN_3414; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3416 = 8'h52 == _T_553 ? 8'h0 : _GEN_3415; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3417 = 8'h53 == _T_553 ? 8'hed : _GEN_3416; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3418 = 8'h54 == _T_553 ? 8'h20 : _GEN_3417; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3419 = 8'h55 == _T_553 ? 8'hfc : _GEN_3418; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3420 = 8'h56 == _T_553 ? 8'hb1 : _GEN_3419; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3421 = 8'h57 == _T_553 ? 8'h5b : _GEN_3420; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3422 = 8'h58 == _T_553 ? 8'h6a : _GEN_3421; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3423 = 8'h59 == _T_553 ? 8'hcb : _GEN_3422; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3424 = 8'h5a == _T_553 ? 8'hbe : _GEN_3423; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3425 = 8'h5b == _T_553 ? 8'h39 : _GEN_3424; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3426 = 8'h5c == _T_553 ? 8'h4a : _GEN_3425; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3427 = 8'h5d == _T_553 ? 8'h4c : _GEN_3426; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3428 = 8'h5e == _T_553 ? 8'h58 : _GEN_3427; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3429 = 8'h5f == _T_553 ? 8'hcf : _GEN_3428; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3430 = 8'h60 == _T_553 ? 8'hd0 : _GEN_3429; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3431 = 8'h61 == _T_553 ? 8'hef : _GEN_3430; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3432 = 8'h62 == _T_553 ? 8'haa : _GEN_3431; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3433 = 8'h63 == _T_553 ? 8'hfb : _GEN_3432; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3434 = 8'h64 == _T_553 ? 8'h43 : _GEN_3433; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3435 = 8'h65 == _T_553 ? 8'h4d : _GEN_3434; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3436 = 8'h66 == _T_553 ? 8'h33 : _GEN_3435; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3437 = 8'h67 == _T_553 ? 8'h85 : _GEN_3436; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3438 = 8'h68 == _T_553 ? 8'h45 : _GEN_3437; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3439 = 8'h69 == _T_553 ? 8'hf9 : _GEN_3438; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3440 = 8'h6a == _T_553 ? 8'h2 : _GEN_3439; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3441 = 8'h6b == _T_553 ? 8'h7f : _GEN_3440; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3442 = 8'h6c == _T_553 ? 8'h50 : _GEN_3441; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3443 = 8'h6d == _T_553 ? 8'h3c : _GEN_3442; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3444 = 8'h6e == _T_553 ? 8'h9f : _GEN_3443; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3445 = 8'h6f == _T_553 ? 8'ha8 : _GEN_3444; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3446 = 8'h70 == _T_553 ? 8'h51 : _GEN_3445; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3447 = 8'h71 == _T_553 ? 8'ha3 : _GEN_3446; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3448 = 8'h72 == _T_553 ? 8'h40 : _GEN_3447; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3449 = 8'h73 == _T_553 ? 8'h8f : _GEN_3448; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3450 = 8'h74 == _T_553 ? 8'h92 : _GEN_3449; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3451 = 8'h75 == _T_553 ? 8'h9d : _GEN_3450; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3452 = 8'h76 == _T_553 ? 8'h38 : _GEN_3451; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3453 = 8'h77 == _T_553 ? 8'hf5 : _GEN_3452; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3454 = 8'h78 == _T_553 ? 8'hbc : _GEN_3453; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3455 = 8'h79 == _T_553 ? 8'hb6 : _GEN_3454; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3456 = 8'h7a == _T_553 ? 8'hda : _GEN_3455; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3457 = 8'h7b == _T_553 ? 8'h21 : _GEN_3456; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3458 = 8'h7c == _T_553 ? 8'h10 : _GEN_3457; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3459 = 8'h7d == _T_553 ? 8'hff : _GEN_3458; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3460 = 8'h7e == _T_553 ? 8'hf3 : _GEN_3459; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3461 = 8'h7f == _T_553 ? 8'hd2 : _GEN_3460; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3462 = 8'h80 == _T_553 ? 8'hcd : _GEN_3461; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3463 = 8'h81 == _T_553 ? 8'hc : _GEN_3462; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3464 = 8'h82 == _T_553 ? 8'h13 : _GEN_3463; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3465 = 8'h83 == _T_553 ? 8'hec : _GEN_3464; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3466 = 8'h84 == _T_553 ? 8'h5f : _GEN_3465; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3467 = 8'h85 == _T_553 ? 8'h97 : _GEN_3466; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3468 = 8'h86 == _T_553 ? 8'h44 : _GEN_3467; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3469 = 8'h87 == _T_553 ? 8'h17 : _GEN_3468; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3470 = 8'h88 == _T_553 ? 8'hc4 : _GEN_3469; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3471 = 8'h89 == _T_553 ? 8'ha7 : _GEN_3470; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3472 = 8'h8a == _T_553 ? 8'h7e : _GEN_3471; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3473 = 8'h8b == _T_553 ? 8'h3d : _GEN_3472; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3474 = 8'h8c == _T_553 ? 8'h64 : _GEN_3473; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3475 = 8'h8d == _T_553 ? 8'h5d : _GEN_3474; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3476 = 8'h8e == _T_553 ? 8'h19 : _GEN_3475; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3477 = 8'h8f == _T_553 ? 8'h73 : _GEN_3476; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3478 = 8'h90 == _T_553 ? 8'h60 : _GEN_3477; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3479 = 8'h91 == _T_553 ? 8'h81 : _GEN_3478; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3480 = 8'h92 == _T_553 ? 8'h4f : _GEN_3479; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3481 = 8'h93 == _T_553 ? 8'hdc : _GEN_3480; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3482 = 8'h94 == _T_553 ? 8'h22 : _GEN_3481; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3483 = 8'h95 == _T_553 ? 8'h2a : _GEN_3482; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3484 = 8'h96 == _T_553 ? 8'h90 : _GEN_3483; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3485 = 8'h97 == _T_553 ? 8'h88 : _GEN_3484; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3486 = 8'h98 == _T_553 ? 8'h46 : _GEN_3485; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3487 = 8'h99 == _T_553 ? 8'hee : _GEN_3486; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3488 = 8'h9a == _T_553 ? 8'hb8 : _GEN_3487; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3489 = 8'h9b == _T_553 ? 8'h14 : _GEN_3488; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3490 = 8'h9c == _T_553 ? 8'hde : _GEN_3489; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3491 = 8'h9d == _T_553 ? 8'h5e : _GEN_3490; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3492 = 8'h9e == _T_553 ? 8'hb : _GEN_3491; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3493 = 8'h9f == _T_553 ? 8'hdb : _GEN_3492; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3494 = 8'ha0 == _T_553 ? 8'he0 : _GEN_3493; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3495 = 8'ha1 == _T_553 ? 8'h32 : _GEN_3494; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3496 = 8'ha2 == _T_553 ? 8'h3a : _GEN_3495; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3497 = 8'ha3 == _T_553 ? 8'ha : _GEN_3496; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3498 = 8'ha4 == _T_553 ? 8'h49 : _GEN_3497; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3499 = 8'ha5 == _T_553 ? 8'h6 : _GEN_3498; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3500 = 8'ha6 == _T_553 ? 8'h24 : _GEN_3499; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3501 = 8'ha7 == _T_553 ? 8'h5c : _GEN_3500; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3502 = 8'ha8 == _T_553 ? 8'hc2 : _GEN_3501; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3503 = 8'ha9 == _T_553 ? 8'hd3 : _GEN_3502; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3504 = 8'haa == _T_553 ? 8'hac : _GEN_3503; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3505 = 8'hab == _T_553 ? 8'h62 : _GEN_3504; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3506 = 8'hac == _T_553 ? 8'h91 : _GEN_3505; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3507 = 8'had == _T_553 ? 8'h95 : _GEN_3506; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3508 = 8'hae == _T_553 ? 8'he4 : _GEN_3507; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3509 = 8'haf == _T_553 ? 8'h79 : _GEN_3508; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3510 = 8'hb0 == _T_553 ? 8'he7 : _GEN_3509; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3511 = 8'hb1 == _T_553 ? 8'hc8 : _GEN_3510; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3512 = 8'hb2 == _T_553 ? 8'h37 : _GEN_3511; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3513 = 8'hb3 == _T_553 ? 8'h6d : _GEN_3512; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3514 = 8'hb4 == _T_553 ? 8'h8d : _GEN_3513; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3515 = 8'hb5 == _T_553 ? 8'hd5 : _GEN_3514; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3516 = 8'hb6 == _T_553 ? 8'h4e : _GEN_3515; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3517 = 8'hb7 == _T_553 ? 8'ha9 : _GEN_3516; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3518 = 8'hb8 == _T_553 ? 8'h6c : _GEN_3517; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3519 = 8'hb9 == _T_553 ? 8'h56 : _GEN_3518; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3520 = 8'hba == _T_553 ? 8'hf4 : _GEN_3519; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3521 = 8'hbb == _T_553 ? 8'hea : _GEN_3520; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3522 = 8'hbc == _T_553 ? 8'h65 : _GEN_3521; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3523 = 8'hbd == _T_553 ? 8'h7a : _GEN_3522; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3524 = 8'hbe == _T_553 ? 8'hae : _GEN_3523; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3525 = 8'hbf == _T_553 ? 8'h8 : _GEN_3524; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3526 = 8'hc0 == _T_553 ? 8'hba : _GEN_3525; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3527 = 8'hc1 == _T_553 ? 8'h78 : _GEN_3526; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3528 = 8'hc2 == _T_553 ? 8'h25 : _GEN_3527; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3529 = 8'hc3 == _T_553 ? 8'h2e : _GEN_3528; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3530 = 8'hc4 == _T_553 ? 8'h1c : _GEN_3529; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3531 = 8'hc5 == _T_553 ? 8'ha6 : _GEN_3530; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3532 = 8'hc6 == _T_553 ? 8'hb4 : _GEN_3531; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3533 = 8'hc7 == _T_553 ? 8'hc6 : _GEN_3532; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3534 = 8'hc8 == _T_553 ? 8'he8 : _GEN_3533; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3535 = 8'hc9 == _T_553 ? 8'hdd : _GEN_3534; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3536 = 8'hca == _T_553 ? 8'h74 : _GEN_3535; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3537 = 8'hcb == _T_553 ? 8'h1f : _GEN_3536; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3538 = 8'hcc == _T_553 ? 8'h4b : _GEN_3537; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3539 = 8'hcd == _T_553 ? 8'hbd : _GEN_3538; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3540 = 8'hce == _T_553 ? 8'h8b : _GEN_3539; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3541 = 8'hcf == _T_553 ? 8'h8a : _GEN_3540; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3542 = 8'hd0 == _T_553 ? 8'h70 : _GEN_3541; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3543 = 8'hd1 == _T_553 ? 8'h3e : _GEN_3542; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3544 = 8'hd2 == _T_553 ? 8'hb5 : _GEN_3543; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3545 = 8'hd3 == _T_553 ? 8'h66 : _GEN_3544; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3546 = 8'hd4 == _T_553 ? 8'h48 : _GEN_3545; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3547 = 8'hd5 == _T_553 ? 8'h3 : _GEN_3546; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3548 = 8'hd6 == _T_553 ? 8'hf6 : _GEN_3547; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3549 = 8'hd7 == _T_553 ? 8'he : _GEN_3548; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3550 = 8'hd8 == _T_553 ? 8'h61 : _GEN_3549; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3551 = 8'hd9 == _T_553 ? 8'h35 : _GEN_3550; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3552 = 8'hda == _T_553 ? 8'h57 : _GEN_3551; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3553 = 8'hdb == _T_553 ? 8'hb9 : _GEN_3552; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3554 = 8'hdc == _T_553 ? 8'h86 : _GEN_3553; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3555 = 8'hdd == _T_553 ? 8'hc1 : _GEN_3554; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3556 = 8'hde == _T_553 ? 8'h1d : _GEN_3555; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3557 = 8'hdf == _T_553 ? 8'h9e : _GEN_3556; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3558 = 8'he0 == _T_553 ? 8'he1 : _GEN_3557; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3559 = 8'he1 == _T_553 ? 8'hf8 : _GEN_3558; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3560 = 8'he2 == _T_553 ? 8'h98 : _GEN_3559; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3561 = 8'he3 == _T_553 ? 8'h11 : _GEN_3560; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3562 = 8'he4 == _T_553 ? 8'h69 : _GEN_3561; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3563 = 8'he5 == _T_553 ? 8'hd9 : _GEN_3562; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3564 = 8'he6 == _T_553 ? 8'h8e : _GEN_3563; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3565 = 8'he7 == _T_553 ? 8'h94 : _GEN_3564; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3566 = 8'he8 == _T_553 ? 8'h9b : _GEN_3565; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3567 = 8'he9 == _T_553 ? 8'h1e : _GEN_3566; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3568 = 8'hea == _T_553 ? 8'h87 : _GEN_3567; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3569 = 8'heb == _T_553 ? 8'he9 : _GEN_3568; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3570 = 8'hec == _T_553 ? 8'hce : _GEN_3569; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3571 = 8'hed == _T_553 ? 8'h55 : _GEN_3570; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3572 = 8'hee == _T_553 ? 8'h28 : _GEN_3571; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3573 = 8'hef == _T_553 ? 8'hdf : _GEN_3572; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3574 = 8'hf0 == _T_553 ? 8'h8c : _GEN_3573; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3575 = 8'hf1 == _T_553 ? 8'ha1 : _GEN_3574; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3576 = 8'hf2 == _T_553 ? 8'h89 : _GEN_3575; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3577 = 8'hf3 == _T_553 ? 8'hd : _GEN_3576; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3578 = 8'hf4 == _T_553 ? 8'hbf : _GEN_3577; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3579 = 8'hf5 == _T_553 ? 8'he6 : _GEN_3578; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3580 = 8'hf6 == _T_553 ? 8'h42 : _GEN_3579; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3581 = 8'hf7 == _T_553 ? 8'h68 : _GEN_3580; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3582 = 8'hf8 == _T_553 ? 8'h41 : _GEN_3581; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3583 = 8'hf9 == _T_553 ? 8'h99 : _GEN_3582; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3584 = 8'hfa == _T_553 ? 8'h2d : _GEN_3583; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3585 = 8'hfb == _T_553 ? 8'hf : _GEN_3584; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3586 = 8'hfc == _T_553 ? 8'hb0 : _GEN_3585; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3587 = 8'hfd == _T_553 ? 8'h54 : _GEN_3586; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3588 = 8'hfe == _T_553 ? 8'hbb : _GEN_3587; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3589 = 8'hff == _T_553 ? 8'h16 : _GEN_3588; // @[Cat.scala 30:58:@2087.4]
  assign _T_561 = {_GEN_3334,_GEN_3589}; // @[Cat.scala 30:58:@2087.4]
  assign _GEN_3590 = 8'h1 == _T_559 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3591 = 8'h2 == _T_559 ? 8'h77 : _GEN_3590; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3592 = 8'h3 == _T_559 ? 8'h7b : _GEN_3591; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3593 = 8'h4 == _T_559 ? 8'hf2 : _GEN_3592; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3594 = 8'h5 == _T_559 ? 8'h6b : _GEN_3593; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3595 = 8'h6 == _T_559 ? 8'h6f : _GEN_3594; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3596 = 8'h7 == _T_559 ? 8'hc5 : _GEN_3595; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3597 = 8'h8 == _T_559 ? 8'h30 : _GEN_3596; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3598 = 8'h9 == _T_559 ? 8'h1 : _GEN_3597; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3599 = 8'ha == _T_559 ? 8'h67 : _GEN_3598; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3600 = 8'hb == _T_559 ? 8'h2b : _GEN_3599; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3601 = 8'hc == _T_559 ? 8'hfe : _GEN_3600; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3602 = 8'hd == _T_559 ? 8'hd7 : _GEN_3601; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3603 = 8'he == _T_559 ? 8'hab : _GEN_3602; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3604 = 8'hf == _T_559 ? 8'h76 : _GEN_3603; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3605 = 8'h10 == _T_559 ? 8'hca : _GEN_3604; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3606 = 8'h11 == _T_559 ? 8'h82 : _GEN_3605; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3607 = 8'h12 == _T_559 ? 8'hc9 : _GEN_3606; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3608 = 8'h13 == _T_559 ? 8'h7d : _GEN_3607; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3609 = 8'h14 == _T_559 ? 8'hfa : _GEN_3608; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3610 = 8'h15 == _T_559 ? 8'h59 : _GEN_3609; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3611 = 8'h16 == _T_559 ? 8'h47 : _GEN_3610; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3612 = 8'h17 == _T_559 ? 8'hf0 : _GEN_3611; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3613 = 8'h18 == _T_559 ? 8'had : _GEN_3612; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3614 = 8'h19 == _T_559 ? 8'hd4 : _GEN_3613; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3615 = 8'h1a == _T_559 ? 8'ha2 : _GEN_3614; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3616 = 8'h1b == _T_559 ? 8'haf : _GEN_3615; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3617 = 8'h1c == _T_559 ? 8'h9c : _GEN_3616; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3618 = 8'h1d == _T_559 ? 8'ha4 : _GEN_3617; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3619 = 8'h1e == _T_559 ? 8'h72 : _GEN_3618; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3620 = 8'h1f == _T_559 ? 8'hc0 : _GEN_3619; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3621 = 8'h20 == _T_559 ? 8'hb7 : _GEN_3620; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3622 = 8'h21 == _T_559 ? 8'hfd : _GEN_3621; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3623 = 8'h22 == _T_559 ? 8'h93 : _GEN_3622; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3624 = 8'h23 == _T_559 ? 8'h26 : _GEN_3623; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3625 = 8'h24 == _T_559 ? 8'h36 : _GEN_3624; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3626 = 8'h25 == _T_559 ? 8'h3f : _GEN_3625; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3627 = 8'h26 == _T_559 ? 8'hf7 : _GEN_3626; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3628 = 8'h27 == _T_559 ? 8'hcc : _GEN_3627; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3629 = 8'h28 == _T_559 ? 8'h34 : _GEN_3628; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3630 = 8'h29 == _T_559 ? 8'ha5 : _GEN_3629; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3631 = 8'h2a == _T_559 ? 8'he5 : _GEN_3630; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3632 = 8'h2b == _T_559 ? 8'hf1 : _GEN_3631; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3633 = 8'h2c == _T_559 ? 8'h71 : _GEN_3632; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3634 = 8'h2d == _T_559 ? 8'hd8 : _GEN_3633; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3635 = 8'h2e == _T_559 ? 8'h31 : _GEN_3634; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3636 = 8'h2f == _T_559 ? 8'h15 : _GEN_3635; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3637 = 8'h30 == _T_559 ? 8'h4 : _GEN_3636; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3638 = 8'h31 == _T_559 ? 8'hc7 : _GEN_3637; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3639 = 8'h32 == _T_559 ? 8'h23 : _GEN_3638; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3640 = 8'h33 == _T_559 ? 8'hc3 : _GEN_3639; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3641 = 8'h34 == _T_559 ? 8'h18 : _GEN_3640; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3642 = 8'h35 == _T_559 ? 8'h96 : _GEN_3641; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3643 = 8'h36 == _T_559 ? 8'h5 : _GEN_3642; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3644 = 8'h37 == _T_559 ? 8'h9a : _GEN_3643; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3645 = 8'h38 == _T_559 ? 8'h7 : _GEN_3644; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3646 = 8'h39 == _T_559 ? 8'h12 : _GEN_3645; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3647 = 8'h3a == _T_559 ? 8'h80 : _GEN_3646; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3648 = 8'h3b == _T_559 ? 8'he2 : _GEN_3647; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3649 = 8'h3c == _T_559 ? 8'heb : _GEN_3648; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3650 = 8'h3d == _T_559 ? 8'h27 : _GEN_3649; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3651 = 8'h3e == _T_559 ? 8'hb2 : _GEN_3650; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3652 = 8'h3f == _T_559 ? 8'h75 : _GEN_3651; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3653 = 8'h40 == _T_559 ? 8'h9 : _GEN_3652; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3654 = 8'h41 == _T_559 ? 8'h83 : _GEN_3653; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3655 = 8'h42 == _T_559 ? 8'h2c : _GEN_3654; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3656 = 8'h43 == _T_559 ? 8'h1a : _GEN_3655; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3657 = 8'h44 == _T_559 ? 8'h1b : _GEN_3656; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3658 = 8'h45 == _T_559 ? 8'h6e : _GEN_3657; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3659 = 8'h46 == _T_559 ? 8'h5a : _GEN_3658; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3660 = 8'h47 == _T_559 ? 8'ha0 : _GEN_3659; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3661 = 8'h48 == _T_559 ? 8'h52 : _GEN_3660; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3662 = 8'h49 == _T_559 ? 8'h3b : _GEN_3661; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3663 = 8'h4a == _T_559 ? 8'hd6 : _GEN_3662; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3664 = 8'h4b == _T_559 ? 8'hb3 : _GEN_3663; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3665 = 8'h4c == _T_559 ? 8'h29 : _GEN_3664; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3666 = 8'h4d == _T_559 ? 8'he3 : _GEN_3665; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3667 = 8'h4e == _T_559 ? 8'h2f : _GEN_3666; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3668 = 8'h4f == _T_559 ? 8'h84 : _GEN_3667; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3669 = 8'h50 == _T_559 ? 8'h53 : _GEN_3668; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3670 = 8'h51 == _T_559 ? 8'hd1 : _GEN_3669; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3671 = 8'h52 == _T_559 ? 8'h0 : _GEN_3670; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3672 = 8'h53 == _T_559 ? 8'hed : _GEN_3671; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3673 = 8'h54 == _T_559 ? 8'h20 : _GEN_3672; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3674 = 8'h55 == _T_559 ? 8'hfc : _GEN_3673; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3675 = 8'h56 == _T_559 ? 8'hb1 : _GEN_3674; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3676 = 8'h57 == _T_559 ? 8'h5b : _GEN_3675; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3677 = 8'h58 == _T_559 ? 8'h6a : _GEN_3676; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3678 = 8'h59 == _T_559 ? 8'hcb : _GEN_3677; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3679 = 8'h5a == _T_559 ? 8'hbe : _GEN_3678; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3680 = 8'h5b == _T_559 ? 8'h39 : _GEN_3679; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3681 = 8'h5c == _T_559 ? 8'h4a : _GEN_3680; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3682 = 8'h5d == _T_559 ? 8'h4c : _GEN_3681; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3683 = 8'h5e == _T_559 ? 8'h58 : _GEN_3682; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3684 = 8'h5f == _T_559 ? 8'hcf : _GEN_3683; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3685 = 8'h60 == _T_559 ? 8'hd0 : _GEN_3684; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3686 = 8'h61 == _T_559 ? 8'hef : _GEN_3685; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3687 = 8'h62 == _T_559 ? 8'haa : _GEN_3686; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3688 = 8'h63 == _T_559 ? 8'hfb : _GEN_3687; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3689 = 8'h64 == _T_559 ? 8'h43 : _GEN_3688; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3690 = 8'h65 == _T_559 ? 8'h4d : _GEN_3689; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3691 = 8'h66 == _T_559 ? 8'h33 : _GEN_3690; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3692 = 8'h67 == _T_559 ? 8'h85 : _GEN_3691; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3693 = 8'h68 == _T_559 ? 8'h45 : _GEN_3692; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3694 = 8'h69 == _T_559 ? 8'hf9 : _GEN_3693; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3695 = 8'h6a == _T_559 ? 8'h2 : _GEN_3694; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3696 = 8'h6b == _T_559 ? 8'h7f : _GEN_3695; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3697 = 8'h6c == _T_559 ? 8'h50 : _GEN_3696; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3698 = 8'h6d == _T_559 ? 8'h3c : _GEN_3697; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3699 = 8'h6e == _T_559 ? 8'h9f : _GEN_3698; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3700 = 8'h6f == _T_559 ? 8'ha8 : _GEN_3699; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3701 = 8'h70 == _T_559 ? 8'h51 : _GEN_3700; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3702 = 8'h71 == _T_559 ? 8'ha3 : _GEN_3701; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3703 = 8'h72 == _T_559 ? 8'h40 : _GEN_3702; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3704 = 8'h73 == _T_559 ? 8'h8f : _GEN_3703; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3705 = 8'h74 == _T_559 ? 8'h92 : _GEN_3704; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3706 = 8'h75 == _T_559 ? 8'h9d : _GEN_3705; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3707 = 8'h76 == _T_559 ? 8'h38 : _GEN_3706; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3708 = 8'h77 == _T_559 ? 8'hf5 : _GEN_3707; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3709 = 8'h78 == _T_559 ? 8'hbc : _GEN_3708; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3710 = 8'h79 == _T_559 ? 8'hb6 : _GEN_3709; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3711 = 8'h7a == _T_559 ? 8'hda : _GEN_3710; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3712 = 8'h7b == _T_559 ? 8'h21 : _GEN_3711; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3713 = 8'h7c == _T_559 ? 8'h10 : _GEN_3712; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3714 = 8'h7d == _T_559 ? 8'hff : _GEN_3713; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3715 = 8'h7e == _T_559 ? 8'hf3 : _GEN_3714; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3716 = 8'h7f == _T_559 ? 8'hd2 : _GEN_3715; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3717 = 8'h80 == _T_559 ? 8'hcd : _GEN_3716; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3718 = 8'h81 == _T_559 ? 8'hc : _GEN_3717; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3719 = 8'h82 == _T_559 ? 8'h13 : _GEN_3718; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3720 = 8'h83 == _T_559 ? 8'hec : _GEN_3719; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3721 = 8'h84 == _T_559 ? 8'h5f : _GEN_3720; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3722 = 8'h85 == _T_559 ? 8'h97 : _GEN_3721; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3723 = 8'h86 == _T_559 ? 8'h44 : _GEN_3722; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3724 = 8'h87 == _T_559 ? 8'h17 : _GEN_3723; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3725 = 8'h88 == _T_559 ? 8'hc4 : _GEN_3724; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3726 = 8'h89 == _T_559 ? 8'ha7 : _GEN_3725; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3727 = 8'h8a == _T_559 ? 8'h7e : _GEN_3726; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3728 = 8'h8b == _T_559 ? 8'h3d : _GEN_3727; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3729 = 8'h8c == _T_559 ? 8'h64 : _GEN_3728; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3730 = 8'h8d == _T_559 ? 8'h5d : _GEN_3729; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3731 = 8'h8e == _T_559 ? 8'h19 : _GEN_3730; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3732 = 8'h8f == _T_559 ? 8'h73 : _GEN_3731; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3733 = 8'h90 == _T_559 ? 8'h60 : _GEN_3732; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3734 = 8'h91 == _T_559 ? 8'h81 : _GEN_3733; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3735 = 8'h92 == _T_559 ? 8'h4f : _GEN_3734; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3736 = 8'h93 == _T_559 ? 8'hdc : _GEN_3735; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3737 = 8'h94 == _T_559 ? 8'h22 : _GEN_3736; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3738 = 8'h95 == _T_559 ? 8'h2a : _GEN_3737; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3739 = 8'h96 == _T_559 ? 8'h90 : _GEN_3738; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3740 = 8'h97 == _T_559 ? 8'h88 : _GEN_3739; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3741 = 8'h98 == _T_559 ? 8'h46 : _GEN_3740; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3742 = 8'h99 == _T_559 ? 8'hee : _GEN_3741; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3743 = 8'h9a == _T_559 ? 8'hb8 : _GEN_3742; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3744 = 8'h9b == _T_559 ? 8'h14 : _GEN_3743; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3745 = 8'h9c == _T_559 ? 8'hde : _GEN_3744; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3746 = 8'h9d == _T_559 ? 8'h5e : _GEN_3745; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3747 = 8'h9e == _T_559 ? 8'hb : _GEN_3746; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3748 = 8'h9f == _T_559 ? 8'hdb : _GEN_3747; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3749 = 8'ha0 == _T_559 ? 8'he0 : _GEN_3748; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3750 = 8'ha1 == _T_559 ? 8'h32 : _GEN_3749; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3751 = 8'ha2 == _T_559 ? 8'h3a : _GEN_3750; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3752 = 8'ha3 == _T_559 ? 8'ha : _GEN_3751; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3753 = 8'ha4 == _T_559 ? 8'h49 : _GEN_3752; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3754 = 8'ha5 == _T_559 ? 8'h6 : _GEN_3753; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3755 = 8'ha6 == _T_559 ? 8'h24 : _GEN_3754; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3756 = 8'ha7 == _T_559 ? 8'h5c : _GEN_3755; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3757 = 8'ha8 == _T_559 ? 8'hc2 : _GEN_3756; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3758 = 8'ha9 == _T_559 ? 8'hd3 : _GEN_3757; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3759 = 8'haa == _T_559 ? 8'hac : _GEN_3758; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3760 = 8'hab == _T_559 ? 8'h62 : _GEN_3759; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3761 = 8'hac == _T_559 ? 8'h91 : _GEN_3760; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3762 = 8'had == _T_559 ? 8'h95 : _GEN_3761; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3763 = 8'hae == _T_559 ? 8'he4 : _GEN_3762; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3764 = 8'haf == _T_559 ? 8'h79 : _GEN_3763; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3765 = 8'hb0 == _T_559 ? 8'he7 : _GEN_3764; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3766 = 8'hb1 == _T_559 ? 8'hc8 : _GEN_3765; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3767 = 8'hb2 == _T_559 ? 8'h37 : _GEN_3766; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3768 = 8'hb3 == _T_559 ? 8'h6d : _GEN_3767; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3769 = 8'hb4 == _T_559 ? 8'h8d : _GEN_3768; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3770 = 8'hb5 == _T_559 ? 8'hd5 : _GEN_3769; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3771 = 8'hb6 == _T_559 ? 8'h4e : _GEN_3770; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3772 = 8'hb7 == _T_559 ? 8'ha9 : _GEN_3771; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3773 = 8'hb8 == _T_559 ? 8'h6c : _GEN_3772; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3774 = 8'hb9 == _T_559 ? 8'h56 : _GEN_3773; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3775 = 8'hba == _T_559 ? 8'hf4 : _GEN_3774; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3776 = 8'hbb == _T_559 ? 8'hea : _GEN_3775; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3777 = 8'hbc == _T_559 ? 8'h65 : _GEN_3776; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3778 = 8'hbd == _T_559 ? 8'h7a : _GEN_3777; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3779 = 8'hbe == _T_559 ? 8'hae : _GEN_3778; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3780 = 8'hbf == _T_559 ? 8'h8 : _GEN_3779; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3781 = 8'hc0 == _T_559 ? 8'hba : _GEN_3780; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3782 = 8'hc1 == _T_559 ? 8'h78 : _GEN_3781; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3783 = 8'hc2 == _T_559 ? 8'h25 : _GEN_3782; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3784 = 8'hc3 == _T_559 ? 8'h2e : _GEN_3783; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3785 = 8'hc4 == _T_559 ? 8'h1c : _GEN_3784; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3786 = 8'hc5 == _T_559 ? 8'ha6 : _GEN_3785; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3787 = 8'hc6 == _T_559 ? 8'hb4 : _GEN_3786; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3788 = 8'hc7 == _T_559 ? 8'hc6 : _GEN_3787; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3789 = 8'hc8 == _T_559 ? 8'he8 : _GEN_3788; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3790 = 8'hc9 == _T_559 ? 8'hdd : _GEN_3789; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3791 = 8'hca == _T_559 ? 8'h74 : _GEN_3790; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3792 = 8'hcb == _T_559 ? 8'h1f : _GEN_3791; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3793 = 8'hcc == _T_559 ? 8'h4b : _GEN_3792; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3794 = 8'hcd == _T_559 ? 8'hbd : _GEN_3793; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3795 = 8'hce == _T_559 ? 8'h8b : _GEN_3794; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3796 = 8'hcf == _T_559 ? 8'h8a : _GEN_3795; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3797 = 8'hd0 == _T_559 ? 8'h70 : _GEN_3796; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3798 = 8'hd1 == _T_559 ? 8'h3e : _GEN_3797; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3799 = 8'hd2 == _T_559 ? 8'hb5 : _GEN_3798; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3800 = 8'hd3 == _T_559 ? 8'h66 : _GEN_3799; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3801 = 8'hd4 == _T_559 ? 8'h48 : _GEN_3800; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3802 = 8'hd5 == _T_559 ? 8'h3 : _GEN_3801; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3803 = 8'hd6 == _T_559 ? 8'hf6 : _GEN_3802; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3804 = 8'hd7 == _T_559 ? 8'he : _GEN_3803; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3805 = 8'hd8 == _T_559 ? 8'h61 : _GEN_3804; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3806 = 8'hd9 == _T_559 ? 8'h35 : _GEN_3805; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3807 = 8'hda == _T_559 ? 8'h57 : _GEN_3806; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3808 = 8'hdb == _T_559 ? 8'hb9 : _GEN_3807; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3809 = 8'hdc == _T_559 ? 8'h86 : _GEN_3808; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3810 = 8'hdd == _T_559 ? 8'hc1 : _GEN_3809; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3811 = 8'hde == _T_559 ? 8'h1d : _GEN_3810; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3812 = 8'hdf == _T_559 ? 8'h9e : _GEN_3811; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3813 = 8'he0 == _T_559 ? 8'he1 : _GEN_3812; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3814 = 8'he1 == _T_559 ? 8'hf8 : _GEN_3813; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3815 = 8'he2 == _T_559 ? 8'h98 : _GEN_3814; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3816 = 8'he3 == _T_559 ? 8'h11 : _GEN_3815; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3817 = 8'he4 == _T_559 ? 8'h69 : _GEN_3816; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3818 = 8'he5 == _T_559 ? 8'hd9 : _GEN_3817; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3819 = 8'he6 == _T_559 ? 8'h8e : _GEN_3818; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3820 = 8'he7 == _T_559 ? 8'h94 : _GEN_3819; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3821 = 8'he8 == _T_559 ? 8'h9b : _GEN_3820; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3822 = 8'he9 == _T_559 ? 8'h1e : _GEN_3821; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3823 = 8'hea == _T_559 ? 8'h87 : _GEN_3822; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3824 = 8'heb == _T_559 ? 8'he9 : _GEN_3823; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3825 = 8'hec == _T_559 ? 8'hce : _GEN_3824; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3826 = 8'hed == _T_559 ? 8'h55 : _GEN_3825; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3827 = 8'hee == _T_559 ? 8'h28 : _GEN_3826; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3828 = 8'hef == _T_559 ? 8'hdf : _GEN_3827; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3829 = 8'hf0 == _T_559 ? 8'h8c : _GEN_3828; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3830 = 8'hf1 == _T_559 ? 8'ha1 : _GEN_3829; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3831 = 8'hf2 == _T_559 ? 8'h89 : _GEN_3830; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3832 = 8'hf3 == _T_559 ? 8'hd : _GEN_3831; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3833 = 8'hf4 == _T_559 ? 8'hbf : _GEN_3832; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3834 = 8'hf5 == _T_559 ? 8'he6 : _GEN_3833; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3835 = 8'hf6 == _T_559 ? 8'h42 : _GEN_3834; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3836 = 8'hf7 == _T_559 ? 8'h68 : _GEN_3835; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3837 = 8'hf8 == _T_559 ? 8'h41 : _GEN_3836; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3838 = 8'hf9 == _T_559 ? 8'h99 : _GEN_3837; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3839 = 8'hfa == _T_559 ? 8'h2d : _GEN_3838; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3840 = 8'hfb == _T_559 ? 8'hf : _GEN_3839; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3841 = 8'hfc == _T_559 ? 8'hb0 : _GEN_3840; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3842 = 8'hfd == _T_559 ? 8'h54 : _GEN_3841; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3843 = 8'hfe == _T_559 ? 8'hbb : _GEN_3842; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3844 = 8'hff == _T_559 ? 8'h16 : _GEN_3843; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3845 = 8'h1 == _T_557 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3846 = 8'h2 == _T_557 ? 8'h77 : _GEN_3845; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3847 = 8'h3 == _T_557 ? 8'h7b : _GEN_3846; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3848 = 8'h4 == _T_557 ? 8'hf2 : _GEN_3847; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3849 = 8'h5 == _T_557 ? 8'h6b : _GEN_3848; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3850 = 8'h6 == _T_557 ? 8'h6f : _GEN_3849; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3851 = 8'h7 == _T_557 ? 8'hc5 : _GEN_3850; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3852 = 8'h8 == _T_557 ? 8'h30 : _GEN_3851; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3853 = 8'h9 == _T_557 ? 8'h1 : _GEN_3852; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3854 = 8'ha == _T_557 ? 8'h67 : _GEN_3853; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3855 = 8'hb == _T_557 ? 8'h2b : _GEN_3854; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3856 = 8'hc == _T_557 ? 8'hfe : _GEN_3855; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3857 = 8'hd == _T_557 ? 8'hd7 : _GEN_3856; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3858 = 8'he == _T_557 ? 8'hab : _GEN_3857; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3859 = 8'hf == _T_557 ? 8'h76 : _GEN_3858; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3860 = 8'h10 == _T_557 ? 8'hca : _GEN_3859; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3861 = 8'h11 == _T_557 ? 8'h82 : _GEN_3860; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3862 = 8'h12 == _T_557 ? 8'hc9 : _GEN_3861; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3863 = 8'h13 == _T_557 ? 8'h7d : _GEN_3862; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3864 = 8'h14 == _T_557 ? 8'hfa : _GEN_3863; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3865 = 8'h15 == _T_557 ? 8'h59 : _GEN_3864; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3866 = 8'h16 == _T_557 ? 8'h47 : _GEN_3865; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3867 = 8'h17 == _T_557 ? 8'hf0 : _GEN_3866; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3868 = 8'h18 == _T_557 ? 8'had : _GEN_3867; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3869 = 8'h19 == _T_557 ? 8'hd4 : _GEN_3868; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3870 = 8'h1a == _T_557 ? 8'ha2 : _GEN_3869; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3871 = 8'h1b == _T_557 ? 8'haf : _GEN_3870; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3872 = 8'h1c == _T_557 ? 8'h9c : _GEN_3871; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3873 = 8'h1d == _T_557 ? 8'ha4 : _GEN_3872; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3874 = 8'h1e == _T_557 ? 8'h72 : _GEN_3873; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3875 = 8'h1f == _T_557 ? 8'hc0 : _GEN_3874; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3876 = 8'h20 == _T_557 ? 8'hb7 : _GEN_3875; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3877 = 8'h21 == _T_557 ? 8'hfd : _GEN_3876; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3878 = 8'h22 == _T_557 ? 8'h93 : _GEN_3877; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3879 = 8'h23 == _T_557 ? 8'h26 : _GEN_3878; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3880 = 8'h24 == _T_557 ? 8'h36 : _GEN_3879; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3881 = 8'h25 == _T_557 ? 8'h3f : _GEN_3880; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3882 = 8'h26 == _T_557 ? 8'hf7 : _GEN_3881; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3883 = 8'h27 == _T_557 ? 8'hcc : _GEN_3882; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3884 = 8'h28 == _T_557 ? 8'h34 : _GEN_3883; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3885 = 8'h29 == _T_557 ? 8'ha5 : _GEN_3884; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3886 = 8'h2a == _T_557 ? 8'he5 : _GEN_3885; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3887 = 8'h2b == _T_557 ? 8'hf1 : _GEN_3886; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3888 = 8'h2c == _T_557 ? 8'h71 : _GEN_3887; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3889 = 8'h2d == _T_557 ? 8'hd8 : _GEN_3888; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3890 = 8'h2e == _T_557 ? 8'h31 : _GEN_3889; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3891 = 8'h2f == _T_557 ? 8'h15 : _GEN_3890; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3892 = 8'h30 == _T_557 ? 8'h4 : _GEN_3891; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3893 = 8'h31 == _T_557 ? 8'hc7 : _GEN_3892; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3894 = 8'h32 == _T_557 ? 8'h23 : _GEN_3893; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3895 = 8'h33 == _T_557 ? 8'hc3 : _GEN_3894; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3896 = 8'h34 == _T_557 ? 8'h18 : _GEN_3895; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3897 = 8'h35 == _T_557 ? 8'h96 : _GEN_3896; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3898 = 8'h36 == _T_557 ? 8'h5 : _GEN_3897; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3899 = 8'h37 == _T_557 ? 8'h9a : _GEN_3898; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3900 = 8'h38 == _T_557 ? 8'h7 : _GEN_3899; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3901 = 8'h39 == _T_557 ? 8'h12 : _GEN_3900; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3902 = 8'h3a == _T_557 ? 8'h80 : _GEN_3901; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3903 = 8'h3b == _T_557 ? 8'he2 : _GEN_3902; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3904 = 8'h3c == _T_557 ? 8'heb : _GEN_3903; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3905 = 8'h3d == _T_557 ? 8'h27 : _GEN_3904; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3906 = 8'h3e == _T_557 ? 8'hb2 : _GEN_3905; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3907 = 8'h3f == _T_557 ? 8'h75 : _GEN_3906; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3908 = 8'h40 == _T_557 ? 8'h9 : _GEN_3907; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3909 = 8'h41 == _T_557 ? 8'h83 : _GEN_3908; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3910 = 8'h42 == _T_557 ? 8'h2c : _GEN_3909; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3911 = 8'h43 == _T_557 ? 8'h1a : _GEN_3910; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3912 = 8'h44 == _T_557 ? 8'h1b : _GEN_3911; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3913 = 8'h45 == _T_557 ? 8'h6e : _GEN_3912; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3914 = 8'h46 == _T_557 ? 8'h5a : _GEN_3913; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3915 = 8'h47 == _T_557 ? 8'ha0 : _GEN_3914; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3916 = 8'h48 == _T_557 ? 8'h52 : _GEN_3915; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3917 = 8'h49 == _T_557 ? 8'h3b : _GEN_3916; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3918 = 8'h4a == _T_557 ? 8'hd6 : _GEN_3917; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3919 = 8'h4b == _T_557 ? 8'hb3 : _GEN_3918; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3920 = 8'h4c == _T_557 ? 8'h29 : _GEN_3919; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3921 = 8'h4d == _T_557 ? 8'he3 : _GEN_3920; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3922 = 8'h4e == _T_557 ? 8'h2f : _GEN_3921; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3923 = 8'h4f == _T_557 ? 8'h84 : _GEN_3922; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3924 = 8'h50 == _T_557 ? 8'h53 : _GEN_3923; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3925 = 8'h51 == _T_557 ? 8'hd1 : _GEN_3924; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3926 = 8'h52 == _T_557 ? 8'h0 : _GEN_3925; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3927 = 8'h53 == _T_557 ? 8'hed : _GEN_3926; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3928 = 8'h54 == _T_557 ? 8'h20 : _GEN_3927; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3929 = 8'h55 == _T_557 ? 8'hfc : _GEN_3928; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3930 = 8'h56 == _T_557 ? 8'hb1 : _GEN_3929; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3931 = 8'h57 == _T_557 ? 8'h5b : _GEN_3930; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3932 = 8'h58 == _T_557 ? 8'h6a : _GEN_3931; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3933 = 8'h59 == _T_557 ? 8'hcb : _GEN_3932; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3934 = 8'h5a == _T_557 ? 8'hbe : _GEN_3933; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3935 = 8'h5b == _T_557 ? 8'h39 : _GEN_3934; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3936 = 8'h5c == _T_557 ? 8'h4a : _GEN_3935; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3937 = 8'h5d == _T_557 ? 8'h4c : _GEN_3936; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3938 = 8'h5e == _T_557 ? 8'h58 : _GEN_3937; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3939 = 8'h5f == _T_557 ? 8'hcf : _GEN_3938; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3940 = 8'h60 == _T_557 ? 8'hd0 : _GEN_3939; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3941 = 8'h61 == _T_557 ? 8'hef : _GEN_3940; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3942 = 8'h62 == _T_557 ? 8'haa : _GEN_3941; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3943 = 8'h63 == _T_557 ? 8'hfb : _GEN_3942; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3944 = 8'h64 == _T_557 ? 8'h43 : _GEN_3943; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3945 = 8'h65 == _T_557 ? 8'h4d : _GEN_3944; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3946 = 8'h66 == _T_557 ? 8'h33 : _GEN_3945; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3947 = 8'h67 == _T_557 ? 8'h85 : _GEN_3946; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3948 = 8'h68 == _T_557 ? 8'h45 : _GEN_3947; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3949 = 8'h69 == _T_557 ? 8'hf9 : _GEN_3948; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3950 = 8'h6a == _T_557 ? 8'h2 : _GEN_3949; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3951 = 8'h6b == _T_557 ? 8'h7f : _GEN_3950; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3952 = 8'h6c == _T_557 ? 8'h50 : _GEN_3951; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3953 = 8'h6d == _T_557 ? 8'h3c : _GEN_3952; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3954 = 8'h6e == _T_557 ? 8'h9f : _GEN_3953; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3955 = 8'h6f == _T_557 ? 8'ha8 : _GEN_3954; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3956 = 8'h70 == _T_557 ? 8'h51 : _GEN_3955; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3957 = 8'h71 == _T_557 ? 8'ha3 : _GEN_3956; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3958 = 8'h72 == _T_557 ? 8'h40 : _GEN_3957; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3959 = 8'h73 == _T_557 ? 8'h8f : _GEN_3958; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3960 = 8'h74 == _T_557 ? 8'h92 : _GEN_3959; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3961 = 8'h75 == _T_557 ? 8'h9d : _GEN_3960; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3962 = 8'h76 == _T_557 ? 8'h38 : _GEN_3961; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3963 = 8'h77 == _T_557 ? 8'hf5 : _GEN_3962; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3964 = 8'h78 == _T_557 ? 8'hbc : _GEN_3963; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3965 = 8'h79 == _T_557 ? 8'hb6 : _GEN_3964; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3966 = 8'h7a == _T_557 ? 8'hda : _GEN_3965; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3967 = 8'h7b == _T_557 ? 8'h21 : _GEN_3966; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3968 = 8'h7c == _T_557 ? 8'h10 : _GEN_3967; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3969 = 8'h7d == _T_557 ? 8'hff : _GEN_3968; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3970 = 8'h7e == _T_557 ? 8'hf3 : _GEN_3969; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3971 = 8'h7f == _T_557 ? 8'hd2 : _GEN_3970; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3972 = 8'h80 == _T_557 ? 8'hcd : _GEN_3971; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3973 = 8'h81 == _T_557 ? 8'hc : _GEN_3972; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3974 = 8'h82 == _T_557 ? 8'h13 : _GEN_3973; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3975 = 8'h83 == _T_557 ? 8'hec : _GEN_3974; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3976 = 8'h84 == _T_557 ? 8'h5f : _GEN_3975; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3977 = 8'h85 == _T_557 ? 8'h97 : _GEN_3976; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3978 = 8'h86 == _T_557 ? 8'h44 : _GEN_3977; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3979 = 8'h87 == _T_557 ? 8'h17 : _GEN_3978; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3980 = 8'h88 == _T_557 ? 8'hc4 : _GEN_3979; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3981 = 8'h89 == _T_557 ? 8'ha7 : _GEN_3980; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3982 = 8'h8a == _T_557 ? 8'h7e : _GEN_3981; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3983 = 8'h8b == _T_557 ? 8'h3d : _GEN_3982; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3984 = 8'h8c == _T_557 ? 8'h64 : _GEN_3983; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3985 = 8'h8d == _T_557 ? 8'h5d : _GEN_3984; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3986 = 8'h8e == _T_557 ? 8'h19 : _GEN_3985; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3987 = 8'h8f == _T_557 ? 8'h73 : _GEN_3986; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3988 = 8'h90 == _T_557 ? 8'h60 : _GEN_3987; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3989 = 8'h91 == _T_557 ? 8'h81 : _GEN_3988; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3990 = 8'h92 == _T_557 ? 8'h4f : _GEN_3989; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3991 = 8'h93 == _T_557 ? 8'hdc : _GEN_3990; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3992 = 8'h94 == _T_557 ? 8'h22 : _GEN_3991; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3993 = 8'h95 == _T_557 ? 8'h2a : _GEN_3992; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3994 = 8'h96 == _T_557 ? 8'h90 : _GEN_3993; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3995 = 8'h97 == _T_557 ? 8'h88 : _GEN_3994; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3996 = 8'h98 == _T_557 ? 8'h46 : _GEN_3995; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3997 = 8'h99 == _T_557 ? 8'hee : _GEN_3996; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3998 = 8'h9a == _T_557 ? 8'hb8 : _GEN_3997; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_3999 = 8'h9b == _T_557 ? 8'h14 : _GEN_3998; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4000 = 8'h9c == _T_557 ? 8'hde : _GEN_3999; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4001 = 8'h9d == _T_557 ? 8'h5e : _GEN_4000; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4002 = 8'h9e == _T_557 ? 8'hb : _GEN_4001; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4003 = 8'h9f == _T_557 ? 8'hdb : _GEN_4002; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4004 = 8'ha0 == _T_557 ? 8'he0 : _GEN_4003; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4005 = 8'ha1 == _T_557 ? 8'h32 : _GEN_4004; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4006 = 8'ha2 == _T_557 ? 8'h3a : _GEN_4005; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4007 = 8'ha3 == _T_557 ? 8'ha : _GEN_4006; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4008 = 8'ha4 == _T_557 ? 8'h49 : _GEN_4007; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4009 = 8'ha5 == _T_557 ? 8'h6 : _GEN_4008; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4010 = 8'ha6 == _T_557 ? 8'h24 : _GEN_4009; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4011 = 8'ha7 == _T_557 ? 8'h5c : _GEN_4010; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4012 = 8'ha8 == _T_557 ? 8'hc2 : _GEN_4011; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4013 = 8'ha9 == _T_557 ? 8'hd3 : _GEN_4012; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4014 = 8'haa == _T_557 ? 8'hac : _GEN_4013; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4015 = 8'hab == _T_557 ? 8'h62 : _GEN_4014; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4016 = 8'hac == _T_557 ? 8'h91 : _GEN_4015; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4017 = 8'had == _T_557 ? 8'h95 : _GEN_4016; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4018 = 8'hae == _T_557 ? 8'he4 : _GEN_4017; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4019 = 8'haf == _T_557 ? 8'h79 : _GEN_4018; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4020 = 8'hb0 == _T_557 ? 8'he7 : _GEN_4019; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4021 = 8'hb1 == _T_557 ? 8'hc8 : _GEN_4020; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4022 = 8'hb2 == _T_557 ? 8'h37 : _GEN_4021; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4023 = 8'hb3 == _T_557 ? 8'h6d : _GEN_4022; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4024 = 8'hb4 == _T_557 ? 8'h8d : _GEN_4023; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4025 = 8'hb5 == _T_557 ? 8'hd5 : _GEN_4024; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4026 = 8'hb6 == _T_557 ? 8'h4e : _GEN_4025; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4027 = 8'hb7 == _T_557 ? 8'ha9 : _GEN_4026; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4028 = 8'hb8 == _T_557 ? 8'h6c : _GEN_4027; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4029 = 8'hb9 == _T_557 ? 8'h56 : _GEN_4028; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4030 = 8'hba == _T_557 ? 8'hf4 : _GEN_4029; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4031 = 8'hbb == _T_557 ? 8'hea : _GEN_4030; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4032 = 8'hbc == _T_557 ? 8'h65 : _GEN_4031; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4033 = 8'hbd == _T_557 ? 8'h7a : _GEN_4032; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4034 = 8'hbe == _T_557 ? 8'hae : _GEN_4033; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4035 = 8'hbf == _T_557 ? 8'h8 : _GEN_4034; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4036 = 8'hc0 == _T_557 ? 8'hba : _GEN_4035; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4037 = 8'hc1 == _T_557 ? 8'h78 : _GEN_4036; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4038 = 8'hc2 == _T_557 ? 8'h25 : _GEN_4037; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4039 = 8'hc3 == _T_557 ? 8'h2e : _GEN_4038; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4040 = 8'hc4 == _T_557 ? 8'h1c : _GEN_4039; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4041 = 8'hc5 == _T_557 ? 8'ha6 : _GEN_4040; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4042 = 8'hc6 == _T_557 ? 8'hb4 : _GEN_4041; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4043 = 8'hc7 == _T_557 ? 8'hc6 : _GEN_4042; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4044 = 8'hc8 == _T_557 ? 8'he8 : _GEN_4043; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4045 = 8'hc9 == _T_557 ? 8'hdd : _GEN_4044; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4046 = 8'hca == _T_557 ? 8'h74 : _GEN_4045; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4047 = 8'hcb == _T_557 ? 8'h1f : _GEN_4046; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4048 = 8'hcc == _T_557 ? 8'h4b : _GEN_4047; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4049 = 8'hcd == _T_557 ? 8'hbd : _GEN_4048; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4050 = 8'hce == _T_557 ? 8'h8b : _GEN_4049; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4051 = 8'hcf == _T_557 ? 8'h8a : _GEN_4050; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4052 = 8'hd0 == _T_557 ? 8'h70 : _GEN_4051; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4053 = 8'hd1 == _T_557 ? 8'h3e : _GEN_4052; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4054 = 8'hd2 == _T_557 ? 8'hb5 : _GEN_4053; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4055 = 8'hd3 == _T_557 ? 8'h66 : _GEN_4054; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4056 = 8'hd4 == _T_557 ? 8'h48 : _GEN_4055; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4057 = 8'hd5 == _T_557 ? 8'h3 : _GEN_4056; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4058 = 8'hd6 == _T_557 ? 8'hf6 : _GEN_4057; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4059 = 8'hd7 == _T_557 ? 8'he : _GEN_4058; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4060 = 8'hd8 == _T_557 ? 8'h61 : _GEN_4059; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4061 = 8'hd9 == _T_557 ? 8'h35 : _GEN_4060; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4062 = 8'hda == _T_557 ? 8'h57 : _GEN_4061; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4063 = 8'hdb == _T_557 ? 8'hb9 : _GEN_4062; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4064 = 8'hdc == _T_557 ? 8'h86 : _GEN_4063; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4065 = 8'hdd == _T_557 ? 8'hc1 : _GEN_4064; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4066 = 8'hde == _T_557 ? 8'h1d : _GEN_4065; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4067 = 8'hdf == _T_557 ? 8'h9e : _GEN_4066; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4068 = 8'he0 == _T_557 ? 8'he1 : _GEN_4067; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4069 = 8'he1 == _T_557 ? 8'hf8 : _GEN_4068; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4070 = 8'he2 == _T_557 ? 8'h98 : _GEN_4069; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4071 = 8'he3 == _T_557 ? 8'h11 : _GEN_4070; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4072 = 8'he4 == _T_557 ? 8'h69 : _GEN_4071; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4073 = 8'he5 == _T_557 ? 8'hd9 : _GEN_4072; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4074 = 8'he6 == _T_557 ? 8'h8e : _GEN_4073; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4075 = 8'he7 == _T_557 ? 8'h94 : _GEN_4074; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4076 = 8'he8 == _T_557 ? 8'h9b : _GEN_4075; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4077 = 8'he9 == _T_557 ? 8'h1e : _GEN_4076; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4078 = 8'hea == _T_557 ? 8'h87 : _GEN_4077; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4079 = 8'heb == _T_557 ? 8'he9 : _GEN_4078; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4080 = 8'hec == _T_557 ? 8'hce : _GEN_4079; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4081 = 8'hed == _T_557 ? 8'h55 : _GEN_4080; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4082 = 8'hee == _T_557 ? 8'h28 : _GEN_4081; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4083 = 8'hef == _T_557 ? 8'hdf : _GEN_4082; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4084 = 8'hf0 == _T_557 ? 8'h8c : _GEN_4083; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4085 = 8'hf1 == _T_557 ? 8'ha1 : _GEN_4084; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4086 = 8'hf2 == _T_557 ? 8'h89 : _GEN_4085; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4087 = 8'hf3 == _T_557 ? 8'hd : _GEN_4086; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4088 = 8'hf4 == _T_557 ? 8'hbf : _GEN_4087; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4089 = 8'hf5 == _T_557 ? 8'he6 : _GEN_4088; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4090 = 8'hf6 == _T_557 ? 8'h42 : _GEN_4089; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4091 = 8'hf7 == _T_557 ? 8'h68 : _GEN_4090; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4092 = 8'hf8 == _T_557 ? 8'h41 : _GEN_4091; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4093 = 8'hf9 == _T_557 ? 8'h99 : _GEN_4092; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4094 = 8'hfa == _T_557 ? 8'h2d : _GEN_4093; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4095 = 8'hfb == _T_557 ? 8'hf : _GEN_4094; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4096 = 8'hfc == _T_557 ? 8'hb0 : _GEN_4095; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4097 = 8'hfd == _T_557 ? 8'h54 : _GEN_4096; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4098 = 8'hfe == _T_557 ? 8'hbb : _GEN_4097; // @[Cat.scala 30:58:@2088.4]
  assign _GEN_4099 = 8'hff == _T_557 ? 8'h16 : _GEN_4098; // @[Cat.scala 30:58:@2088.4]
  assign _T_562 = {_GEN_3844,_GEN_4099}; // @[Cat.scala 30:58:@2088.4]
  assign x3 = {_T_562,_T_561}; // @[Cat.scala 30:58:@2089.4]
  assign _T_563 = io_addr2[103:96]; // @[sbox.scala 76:26:@2090.4]
  assign _T_565 = io_addr2[111:104]; // @[sbox.scala 77:26:@2091.4]
  assign _T_567 = io_addr2[119:112]; // @[sbox.scala 78:26:@2092.4]
  assign _T_569 = io_addr2[127:120]; // @[sbox.scala 79:26:@2093.4]
  assign _GEN_4100 = 8'h1 == _T_565 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4101 = 8'h2 == _T_565 ? 8'h77 : _GEN_4100; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4102 = 8'h3 == _T_565 ? 8'h7b : _GEN_4101; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4103 = 8'h4 == _T_565 ? 8'hf2 : _GEN_4102; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4104 = 8'h5 == _T_565 ? 8'h6b : _GEN_4103; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4105 = 8'h6 == _T_565 ? 8'h6f : _GEN_4104; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4106 = 8'h7 == _T_565 ? 8'hc5 : _GEN_4105; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4107 = 8'h8 == _T_565 ? 8'h30 : _GEN_4106; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4108 = 8'h9 == _T_565 ? 8'h1 : _GEN_4107; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4109 = 8'ha == _T_565 ? 8'h67 : _GEN_4108; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4110 = 8'hb == _T_565 ? 8'h2b : _GEN_4109; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4111 = 8'hc == _T_565 ? 8'hfe : _GEN_4110; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4112 = 8'hd == _T_565 ? 8'hd7 : _GEN_4111; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4113 = 8'he == _T_565 ? 8'hab : _GEN_4112; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4114 = 8'hf == _T_565 ? 8'h76 : _GEN_4113; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4115 = 8'h10 == _T_565 ? 8'hca : _GEN_4114; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4116 = 8'h11 == _T_565 ? 8'h82 : _GEN_4115; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4117 = 8'h12 == _T_565 ? 8'hc9 : _GEN_4116; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4118 = 8'h13 == _T_565 ? 8'h7d : _GEN_4117; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4119 = 8'h14 == _T_565 ? 8'hfa : _GEN_4118; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4120 = 8'h15 == _T_565 ? 8'h59 : _GEN_4119; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4121 = 8'h16 == _T_565 ? 8'h47 : _GEN_4120; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4122 = 8'h17 == _T_565 ? 8'hf0 : _GEN_4121; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4123 = 8'h18 == _T_565 ? 8'had : _GEN_4122; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4124 = 8'h19 == _T_565 ? 8'hd4 : _GEN_4123; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4125 = 8'h1a == _T_565 ? 8'ha2 : _GEN_4124; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4126 = 8'h1b == _T_565 ? 8'haf : _GEN_4125; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4127 = 8'h1c == _T_565 ? 8'h9c : _GEN_4126; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4128 = 8'h1d == _T_565 ? 8'ha4 : _GEN_4127; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4129 = 8'h1e == _T_565 ? 8'h72 : _GEN_4128; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4130 = 8'h1f == _T_565 ? 8'hc0 : _GEN_4129; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4131 = 8'h20 == _T_565 ? 8'hb7 : _GEN_4130; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4132 = 8'h21 == _T_565 ? 8'hfd : _GEN_4131; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4133 = 8'h22 == _T_565 ? 8'h93 : _GEN_4132; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4134 = 8'h23 == _T_565 ? 8'h26 : _GEN_4133; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4135 = 8'h24 == _T_565 ? 8'h36 : _GEN_4134; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4136 = 8'h25 == _T_565 ? 8'h3f : _GEN_4135; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4137 = 8'h26 == _T_565 ? 8'hf7 : _GEN_4136; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4138 = 8'h27 == _T_565 ? 8'hcc : _GEN_4137; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4139 = 8'h28 == _T_565 ? 8'h34 : _GEN_4138; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4140 = 8'h29 == _T_565 ? 8'ha5 : _GEN_4139; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4141 = 8'h2a == _T_565 ? 8'he5 : _GEN_4140; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4142 = 8'h2b == _T_565 ? 8'hf1 : _GEN_4141; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4143 = 8'h2c == _T_565 ? 8'h71 : _GEN_4142; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4144 = 8'h2d == _T_565 ? 8'hd8 : _GEN_4143; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4145 = 8'h2e == _T_565 ? 8'h31 : _GEN_4144; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4146 = 8'h2f == _T_565 ? 8'h15 : _GEN_4145; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4147 = 8'h30 == _T_565 ? 8'h4 : _GEN_4146; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4148 = 8'h31 == _T_565 ? 8'hc7 : _GEN_4147; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4149 = 8'h32 == _T_565 ? 8'h23 : _GEN_4148; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4150 = 8'h33 == _T_565 ? 8'hc3 : _GEN_4149; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4151 = 8'h34 == _T_565 ? 8'h18 : _GEN_4150; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4152 = 8'h35 == _T_565 ? 8'h96 : _GEN_4151; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4153 = 8'h36 == _T_565 ? 8'h5 : _GEN_4152; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4154 = 8'h37 == _T_565 ? 8'h9a : _GEN_4153; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4155 = 8'h38 == _T_565 ? 8'h7 : _GEN_4154; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4156 = 8'h39 == _T_565 ? 8'h12 : _GEN_4155; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4157 = 8'h3a == _T_565 ? 8'h80 : _GEN_4156; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4158 = 8'h3b == _T_565 ? 8'he2 : _GEN_4157; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4159 = 8'h3c == _T_565 ? 8'heb : _GEN_4158; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4160 = 8'h3d == _T_565 ? 8'h27 : _GEN_4159; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4161 = 8'h3e == _T_565 ? 8'hb2 : _GEN_4160; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4162 = 8'h3f == _T_565 ? 8'h75 : _GEN_4161; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4163 = 8'h40 == _T_565 ? 8'h9 : _GEN_4162; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4164 = 8'h41 == _T_565 ? 8'h83 : _GEN_4163; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4165 = 8'h42 == _T_565 ? 8'h2c : _GEN_4164; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4166 = 8'h43 == _T_565 ? 8'h1a : _GEN_4165; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4167 = 8'h44 == _T_565 ? 8'h1b : _GEN_4166; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4168 = 8'h45 == _T_565 ? 8'h6e : _GEN_4167; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4169 = 8'h46 == _T_565 ? 8'h5a : _GEN_4168; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4170 = 8'h47 == _T_565 ? 8'ha0 : _GEN_4169; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4171 = 8'h48 == _T_565 ? 8'h52 : _GEN_4170; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4172 = 8'h49 == _T_565 ? 8'h3b : _GEN_4171; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4173 = 8'h4a == _T_565 ? 8'hd6 : _GEN_4172; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4174 = 8'h4b == _T_565 ? 8'hb3 : _GEN_4173; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4175 = 8'h4c == _T_565 ? 8'h29 : _GEN_4174; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4176 = 8'h4d == _T_565 ? 8'he3 : _GEN_4175; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4177 = 8'h4e == _T_565 ? 8'h2f : _GEN_4176; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4178 = 8'h4f == _T_565 ? 8'h84 : _GEN_4177; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4179 = 8'h50 == _T_565 ? 8'h53 : _GEN_4178; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4180 = 8'h51 == _T_565 ? 8'hd1 : _GEN_4179; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4181 = 8'h52 == _T_565 ? 8'h0 : _GEN_4180; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4182 = 8'h53 == _T_565 ? 8'hed : _GEN_4181; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4183 = 8'h54 == _T_565 ? 8'h20 : _GEN_4182; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4184 = 8'h55 == _T_565 ? 8'hfc : _GEN_4183; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4185 = 8'h56 == _T_565 ? 8'hb1 : _GEN_4184; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4186 = 8'h57 == _T_565 ? 8'h5b : _GEN_4185; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4187 = 8'h58 == _T_565 ? 8'h6a : _GEN_4186; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4188 = 8'h59 == _T_565 ? 8'hcb : _GEN_4187; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4189 = 8'h5a == _T_565 ? 8'hbe : _GEN_4188; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4190 = 8'h5b == _T_565 ? 8'h39 : _GEN_4189; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4191 = 8'h5c == _T_565 ? 8'h4a : _GEN_4190; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4192 = 8'h5d == _T_565 ? 8'h4c : _GEN_4191; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4193 = 8'h5e == _T_565 ? 8'h58 : _GEN_4192; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4194 = 8'h5f == _T_565 ? 8'hcf : _GEN_4193; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4195 = 8'h60 == _T_565 ? 8'hd0 : _GEN_4194; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4196 = 8'h61 == _T_565 ? 8'hef : _GEN_4195; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4197 = 8'h62 == _T_565 ? 8'haa : _GEN_4196; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4198 = 8'h63 == _T_565 ? 8'hfb : _GEN_4197; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4199 = 8'h64 == _T_565 ? 8'h43 : _GEN_4198; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4200 = 8'h65 == _T_565 ? 8'h4d : _GEN_4199; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4201 = 8'h66 == _T_565 ? 8'h33 : _GEN_4200; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4202 = 8'h67 == _T_565 ? 8'h85 : _GEN_4201; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4203 = 8'h68 == _T_565 ? 8'h45 : _GEN_4202; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4204 = 8'h69 == _T_565 ? 8'hf9 : _GEN_4203; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4205 = 8'h6a == _T_565 ? 8'h2 : _GEN_4204; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4206 = 8'h6b == _T_565 ? 8'h7f : _GEN_4205; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4207 = 8'h6c == _T_565 ? 8'h50 : _GEN_4206; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4208 = 8'h6d == _T_565 ? 8'h3c : _GEN_4207; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4209 = 8'h6e == _T_565 ? 8'h9f : _GEN_4208; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4210 = 8'h6f == _T_565 ? 8'ha8 : _GEN_4209; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4211 = 8'h70 == _T_565 ? 8'h51 : _GEN_4210; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4212 = 8'h71 == _T_565 ? 8'ha3 : _GEN_4211; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4213 = 8'h72 == _T_565 ? 8'h40 : _GEN_4212; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4214 = 8'h73 == _T_565 ? 8'h8f : _GEN_4213; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4215 = 8'h74 == _T_565 ? 8'h92 : _GEN_4214; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4216 = 8'h75 == _T_565 ? 8'h9d : _GEN_4215; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4217 = 8'h76 == _T_565 ? 8'h38 : _GEN_4216; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4218 = 8'h77 == _T_565 ? 8'hf5 : _GEN_4217; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4219 = 8'h78 == _T_565 ? 8'hbc : _GEN_4218; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4220 = 8'h79 == _T_565 ? 8'hb6 : _GEN_4219; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4221 = 8'h7a == _T_565 ? 8'hda : _GEN_4220; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4222 = 8'h7b == _T_565 ? 8'h21 : _GEN_4221; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4223 = 8'h7c == _T_565 ? 8'h10 : _GEN_4222; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4224 = 8'h7d == _T_565 ? 8'hff : _GEN_4223; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4225 = 8'h7e == _T_565 ? 8'hf3 : _GEN_4224; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4226 = 8'h7f == _T_565 ? 8'hd2 : _GEN_4225; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4227 = 8'h80 == _T_565 ? 8'hcd : _GEN_4226; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4228 = 8'h81 == _T_565 ? 8'hc : _GEN_4227; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4229 = 8'h82 == _T_565 ? 8'h13 : _GEN_4228; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4230 = 8'h83 == _T_565 ? 8'hec : _GEN_4229; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4231 = 8'h84 == _T_565 ? 8'h5f : _GEN_4230; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4232 = 8'h85 == _T_565 ? 8'h97 : _GEN_4231; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4233 = 8'h86 == _T_565 ? 8'h44 : _GEN_4232; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4234 = 8'h87 == _T_565 ? 8'h17 : _GEN_4233; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4235 = 8'h88 == _T_565 ? 8'hc4 : _GEN_4234; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4236 = 8'h89 == _T_565 ? 8'ha7 : _GEN_4235; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4237 = 8'h8a == _T_565 ? 8'h7e : _GEN_4236; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4238 = 8'h8b == _T_565 ? 8'h3d : _GEN_4237; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4239 = 8'h8c == _T_565 ? 8'h64 : _GEN_4238; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4240 = 8'h8d == _T_565 ? 8'h5d : _GEN_4239; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4241 = 8'h8e == _T_565 ? 8'h19 : _GEN_4240; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4242 = 8'h8f == _T_565 ? 8'h73 : _GEN_4241; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4243 = 8'h90 == _T_565 ? 8'h60 : _GEN_4242; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4244 = 8'h91 == _T_565 ? 8'h81 : _GEN_4243; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4245 = 8'h92 == _T_565 ? 8'h4f : _GEN_4244; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4246 = 8'h93 == _T_565 ? 8'hdc : _GEN_4245; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4247 = 8'h94 == _T_565 ? 8'h22 : _GEN_4246; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4248 = 8'h95 == _T_565 ? 8'h2a : _GEN_4247; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4249 = 8'h96 == _T_565 ? 8'h90 : _GEN_4248; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4250 = 8'h97 == _T_565 ? 8'h88 : _GEN_4249; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4251 = 8'h98 == _T_565 ? 8'h46 : _GEN_4250; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4252 = 8'h99 == _T_565 ? 8'hee : _GEN_4251; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4253 = 8'h9a == _T_565 ? 8'hb8 : _GEN_4252; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4254 = 8'h9b == _T_565 ? 8'h14 : _GEN_4253; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4255 = 8'h9c == _T_565 ? 8'hde : _GEN_4254; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4256 = 8'h9d == _T_565 ? 8'h5e : _GEN_4255; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4257 = 8'h9e == _T_565 ? 8'hb : _GEN_4256; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4258 = 8'h9f == _T_565 ? 8'hdb : _GEN_4257; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4259 = 8'ha0 == _T_565 ? 8'he0 : _GEN_4258; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4260 = 8'ha1 == _T_565 ? 8'h32 : _GEN_4259; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4261 = 8'ha2 == _T_565 ? 8'h3a : _GEN_4260; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4262 = 8'ha3 == _T_565 ? 8'ha : _GEN_4261; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4263 = 8'ha4 == _T_565 ? 8'h49 : _GEN_4262; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4264 = 8'ha5 == _T_565 ? 8'h6 : _GEN_4263; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4265 = 8'ha6 == _T_565 ? 8'h24 : _GEN_4264; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4266 = 8'ha7 == _T_565 ? 8'h5c : _GEN_4265; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4267 = 8'ha8 == _T_565 ? 8'hc2 : _GEN_4266; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4268 = 8'ha9 == _T_565 ? 8'hd3 : _GEN_4267; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4269 = 8'haa == _T_565 ? 8'hac : _GEN_4268; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4270 = 8'hab == _T_565 ? 8'h62 : _GEN_4269; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4271 = 8'hac == _T_565 ? 8'h91 : _GEN_4270; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4272 = 8'had == _T_565 ? 8'h95 : _GEN_4271; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4273 = 8'hae == _T_565 ? 8'he4 : _GEN_4272; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4274 = 8'haf == _T_565 ? 8'h79 : _GEN_4273; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4275 = 8'hb0 == _T_565 ? 8'he7 : _GEN_4274; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4276 = 8'hb1 == _T_565 ? 8'hc8 : _GEN_4275; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4277 = 8'hb2 == _T_565 ? 8'h37 : _GEN_4276; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4278 = 8'hb3 == _T_565 ? 8'h6d : _GEN_4277; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4279 = 8'hb4 == _T_565 ? 8'h8d : _GEN_4278; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4280 = 8'hb5 == _T_565 ? 8'hd5 : _GEN_4279; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4281 = 8'hb6 == _T_565 ? 8'h4e : _GEN_4280; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4282 = 8'hb7 == _T_565 ? 8'ha9 : _GEN_4281; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4283 = 8'hb8 == _T_565 ? 8'h6c : _GEN_4282; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4284 = 8'hb9 == _T_565 ? 8'h56 : _GEN_4283; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4285 = 8'hba == _T_565 ? 8'hf4 : _GEN_4284; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4286 = 8'hbb == _T_565 ? 8'hea : _GEN_4285; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4287 = 8'hbc == _T_565 ? 8'h65 : _GEN_4286; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4288 = 8'hbd == _T_565 ? 8'h7a : _GEN_4287; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4289 = 8'hbe == _T_565 ? 8'hae : _GEN_4288; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4290 = 8'hbf == _T_565 ? 8'h8 : _GEN_4289; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4291 = 8'hc0 == _T_565 ? 8'hba : _GEN_4290; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4292 = 8'hc1 == _T_565 ? 8'h78 : _GEN_4291; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4293 = 8'hc2 == _T_565 ? 8'h25 : _GEN_4292; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4294 = 8'hc3 == _T_565 ? 8'h2e : _GEN_4293; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4295 = 8'hc4 == _T_565 ? 8'h1c : _GEN_4294; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4296 = 8'hc5 == _T_565 ? 8'ha6 : _GEN_4295; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4297 = 8'hc6 == _T_565 ? 8'hb4 : _GEN_4296; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4298 = 8'hc7 == _T_565 ? 8'hc6 : _GEN_4297; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4299 = 8'hc8 == _T_565 ? 8'he8 : _GEN_4298; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4300 = 8'hc9 == _T_565 ? 8'hdd : _GEN_4299; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4301 = 8'hca == _T_565 ? 8'h74 : _GEN_4300; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4302 = 8'hcb == _T_565 ? 8'h1f : _GEN_4301; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4303 = 8'hcc == _T_565 ? 8'h4b : _GEN_4302; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4304 = 8'hcd == _T_565 ? 8'hbd : _GEN_4303; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4305 = 8'hce == _T_565 ? 8'h8b : _GEN_4304; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4306 = 8'hcf == _T_565 ? 8'h8a : _GEN_4305; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4307 = 8'hd0 == _T_565 ? 8'h70 : _GEN_4306; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4308 = 8'hd1 == _T_565 ? 8'h3e : _GEN_4307; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4309 = 8'hd2 == _T_565 ? 8'hb5 : _GEN_4308; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4310 = 8'hd3 == _T_565 ? 8'h66 : _GEN_4309; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4311 = 8'hd4 == _T_565 ? 8'h48 : _GEN_4310; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4312 = 8'hd5 == _T_565 ? 8'h3 : _GEN_4311; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4313 = 8'hd6 == _T_565 ? 8'hf6 : _GEN_4312; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4314 = 8'hd7 == _T_565 ? 8'he : _GEN_4313; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4315 = 8'hd8 == _T_565 ? 8'h61 : _GEN_4314; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4316 = 8'hd9 == _T_565 ? 8'h35 : _GEN_4315; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4317 = 8'hda == _T_565 ? 8'h57 : _GEN_4316; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4318 = 8'hdb == _T_565 ? 8'hb9 : _GEN_4317; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4319 = 8'hdc == _T_565 ? 8'h86 : _GEN_4318; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4320 = 8'hdd == _T_565 ? 8'hc1 : _GEN_4319; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4321 = 8'hde == _T_565 ? 8'h1d : _GEN_4320; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4322 = 8'hdf == _T_565 ? 8'h9e : _GEN_4321; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4323 = 8'he0 == _T_565 ? 8'he1 : _GEN_4322; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4324 = 8'he1 == _T_565 ? 8'hf8 : _GEN_4323; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4325 = 8'he2 == _T_565 ? 8'h98 : _GEN_4324; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4326 = 8'he3 == _T_565 ? 8'h11 : _GEN_4325; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4327 = 8'he4 == _T_565 ? 8'h69 : _GEN_4326; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4328 = 8'he5 == _T_565 ? 8'hd9 : _GEN_4327; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4329 = 8'he6 == _T_565 ? 8'h8e : _GEN_4328; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4330 = 8'he7 == _T_565 ? 8'h94 : _GEN_4329; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4331 = 8'he8 == _T_565 ? 8'h9b : _GEN_4330; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4332 = 8'he9 == _T_565 ? 8'h1e : _GEN_4331; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4333 = 8'hea == _T_565 ? 8'h87 : _GEN_4332; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4334 = 8'heb == _T_565 ? 8'he9 : _GEN_4333; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4335 = 8'hec == _T_565 ? 8'hce : _GEN_4334; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4336 = 8'hed == _T_565 ? 8'h55 : _GEN_4335; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4337 = 8'hee == _T_565 ? 8'h28 : _GEN_4336; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4338 = 8'hef == _T_565 ? 8'hdf : _GEN_4337; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4339 = 8'hf0 == _T_565 ? 8'h8c : _GEN_4338; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4340 = 8'hf1 == _T_565 ? 8'ha1 : _GEN_4339; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4341 = 8'hf2 == _T_565 ? 8'h89 : _GEN_4340; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4342 = 8'hf3 == _T_565 ? 8'hd : _GEN_4341; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4343 = 8'hf4 == _T_565 ? 8'hbf : _GEN_4342; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4344 = 8'hf5 == _T_565 ? 8'he6 : _GEN_4343; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4345 = 8'hf6 == _T_565 ? 8'h42 : _GEN_4344; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4346 = 8'hf7 == _T_565 ? 8'h68 : _GEN_4345; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4347 = 8'hf8 == _T_565 ? 8'h41 : _GEN_4346; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4348 = 8'hf9 == _T_565 ? 8'h99 : _GEN_4347; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4349 = 8'hfa == _T_565 ? 8'h2d : _GEN_4348; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4350 = 8'hfb == _T_565 ? 8'hf : _GEN_4349; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4351 = 8'hfc == _T_565 ? 8'hb0 : _GEN_4350; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4352 = 8'hfd == _T_565 ? 8'h54 : _GEN_4351; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4353 = 8'hfe == _T_565 ? 8'hbb : _GEN_4352; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4354 = 8'hff == _T_565 ? 8'h16 : _GEN_4353; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4355 = 8'h1 == _T_563 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4356 = 8'h2 == _T_563 ? 8'h77 : _GEN_4355; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4357 = 8'h3 == _T_563 ? 8'h7b : _GEN_4356; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4358 = 8'h4 == _T_563 ? 8'hf2 : _GEN_4357; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4359 = 8'h5 == _T_563 ? 8'h6b : _GEN_4358; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4360 = 8'h6 == _T_563 ? 8'h6f : _GEN_4359; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4361 = 8'h7 == _T_563 ? 8'hc5 : _GEN_4360; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4362 = 8'h8 == _T_563 ? 8'h30 : _GEN_4361; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4363 = 8'h9 == _T_563 ? 8'h1 : _GEN_4362; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4364 = 8'ha == _T_563 ? 8'h67 : _GEN_4363; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4365 = 8'hb == _T_563 ? 8'h2b : _GEN_4364; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4366 = 8'hc == _T_563 ? 8'hfe : _GEN_4365; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4367 = 8'hd == _T_563 ? 8'hd7 : _GEN_4366; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4368 = 8'he == _T_563 ? 8'hab : _GEN_4367; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4369 = 8'hf == _T_563 ? 8'h76 : _GEN_4368; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4370 = 8'h10 == _T_563 ? 8'hca : _GEN_4369; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4371 = 8'h11 == _T_563 ? 8'h82 : _GEN_4370; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4372 = 8'h12 == _T_563 ? 8'hc9 : _GEN_4371; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4373 = 8'h13 == _T_563 ? 8'h7d : _GEN_4372; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4374 = 8'h14 == _T_563 ? 8'hfa : _GEN_4373; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4375 = 8'h15 == _T_563 ? 8'h59 : _GEN_4374; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4376 = 8'h16 == _T_563 ? 8'h47 : _GEN_4375; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4377 = 8'h17 == _T_563 ? 8'hf0 : _GEN_4376; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4378 = 8'h18 == _T_563 ? 8'had : _GEN_4377; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4379 = 8'h19 == _T_563 ? 8'hd4 : _GEN_4378; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4380 = 8'h1a == _T_563 ? 8'ha2 : _GEN_4379; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4381 = 8'h1b == _T_563 ? 8'haf : _GEN_4380; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4382 = 8'h1c == _T_563 ? 8'h9c : _GEN_4381; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4383 = 8'h1d == _T_563 ? 8'ha4 : _GEN_4382; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4384 = 8'h1e == _T_563 ? 8'h72 : _GEN_4383; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4385 = 8'h1f == _T_563 ? 8'hc0 : _GEN_4384; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4386 = 8'h20 == _T_563 ? 8'hb7 : _GEN_4385; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4387 = 8'h21 == _T_563 ? 8'hfd : _GEN_4386; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4388 = 8'h22 == _T_563 ? 8'h93 : _GEN_4387; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4389 = 8'h23 == _T_563 ? 8'h26 : _GEN_4388; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4390 = 8'h24 == _T_563 ? 8'h36 : _GEN_4389; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4391 = 8'h25 == _T_563 ? 8'h3f : _GEN_4390; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4392 = 8'h26 == _T_563 ? 8'hf7 : _GEN_4391; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4393 = 8'h27 == _T_563 ? 8'hcc : _GEN_4392; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4394 = 8'h28 == _T_563 ? 8'h34 : _GEN_4393; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4395 = 8'h29 == _T_563 ? 8'ha5 : _GEN_4394; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4396 = 8'h2a == _T_563 ? 8'he5 : _GEN_4395; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4397 = 8'h2b == _T_563 ? 8'hf1 : _GEN_4396; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4398 = 8'h2c == _T_563 ? 8'h71 : _GEN_4397; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4399 = 8'h2d == _T_563 ? 8'hd8 : _GEN_4398; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4400 = 8'h2e == _T_563 ? 8'h31 : _GEN_4399; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4401 = 8'h2f == _T_563 ? 8'h15 : _GEN_4400; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4402 = 8'h30 == _T_563 ? 8'h4 : _GEN_4401; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4403 = 8'h31 == _T_563 ? 8'hc7 : _GEN_4402; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4404 = 8'h32 == _T_563 ? 8'h23 : _GEN_4403; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4405 = 8'h33 == _T_563 ? 8'hc3 : _GEN_4404; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4406 = 8'h34 == _T_563 ? 8'h18 : _GEN_4405; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4407 = 8'h35 == _T_563 ? 8'h96 : _GEN_4406; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4408 = 8'h36 == _T_563 ? 8'h5 : _GEN_4407; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4409 = 8'h37 == _T_563 ? 8'h9a : _GEN_4408; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4410 = 8'h38 == _T_563 ? 8'h7 : _GEN_4409; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4411 = 8'h39 == _T_563 ? 8'h12 : _GEN_4410; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4412 = 8'h3a == _T_563 ? 8'h80 : _GEN_4411; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4413 = 8'h3b == _T_563 ? 8'he2 : _GEN_4412; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4414 = 8'h3c == _T_563 ? 8'heb : _GEN_4413; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4415 = 8'h3d == _T_563 ? 8'h27 : _GEN_4414; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4416 = 8'h3e == _T_563 ? 8'hb2 : _GEN_4415; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4417 = 8'h3f == _T_563 ? 8'h75 : _GEN_4416; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4418 = 8'h40 == _T_563 ? 8'h9 : _GEN_4417; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4419 = 8'h41 == _T_563 ? 8'h83 : _GEN_4418; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4420 = 8'h42 == _T_563 ? 8'h2c : _GEN_4419; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4421 = 8'h43 == _T_563 ? 8'h1a : _GEN_4420; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4422 = 8'h44 == _T_563 ? 8'h1b : _GEN_4421; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4423 = 8'h45 == _T_563 ? 8'h6e : _GEN_4422; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4424 = 8'h46 == _T_563 ? 8'h5a : _GEN_4423; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4425 = 8'h47 == _T_563 ? 8'ha0 : _GEN_4424; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4426 = 8'h48 == _T_563 ? 8'h52 : _GEN_4425; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4427 = 8'h49 == _T_563 ? 8'h3b : _GEN_4426; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4428 = 8'h4a == _T_563 ? 8'hd6 : _GEN_4427; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4429 = 8'h4b == _T_563 ? 8'hb3 : _GEN_4428; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4430 = 8'h4c == _T_563 ? 8'h29 : _GEN_4429; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4431 = 8'h4d == _T_563 ? 8'he3 : _GEN_4430; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4432 = 8'h4e == _T_563 ? 8'h2f : _GEN_4431; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4433 = 8'h4f == _T_563 ? 8'h84 : _GEN_4432; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4434 = 8'h50 == _T_563 ? 8'h53 : _GEN_4433; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4435 = 8'h51 == _T_563 ? 8'hd1 : _GEN_4434; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4436 = 8'h52 == _T_563 ? 8'h0 : _GEN_4435; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4437 = 8'h53 == _T_563 ? 8'hed : _GEN_4436; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4438 = 8'h54 == _T_563 ? 8'h20 : _GEN_4437; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4439 = 8'h55 == _T_563 ? 8'hfc : _GEN_4438; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4440 = 8'h56 == _T_563 ? 8'hb1 : _GEN_4439; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4441 = 8'h57 == _T_563 ? 8'h5b : _GEN_4440; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4442 = 8'h58 == _T_563 ? 8'h6a : _GEN_4441; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4443 = 8'h59 == _T_563 ? 8'hcb : _GEN_4442; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4444 = 8'h5a == _T_563 ? 8'hbe : _GEN_4443; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4445 = 8'h5b == _T_563 ? 8'h39 : _GEN_4444; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4446 = 8'h5c == _T_563 ? 8'h4a : _GEN_4445; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4447 = 8'h5d == _T_563 ? 8'h4c : _GEN_4446; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4448 = 8'h5e == _T_563 ? 8'h58 : _GEN_4447; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4449 = 8'h5f == _T_563 ? 8'hcf : _GEN_4448; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4450 = 8'h60 == _T_563 ? 8'hd0 : _GEN_4449; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4451 = 8'h61 == _T_563 ? 8'hef : _GEN_4450; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4452 = 8'h62 == _T_563 ? 8'haa : _GEN_4451; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4453 = 8'h63 == _T_563 ? 8'hfb : _GEN_4452; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4454 = 8'h64 == _T_563 ? 8'h43 : _GEN_4453; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4455 = 8'h65 == _T_563 ? 8'h4d : _GEN_4454; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4456 = 8'h66 == _T_563 ? 8'h33 : _GEN_4455; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4457 = 8'h67 == _T_563 ? 8'h85 : _GEN_4456; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4458 = 8'h68 == _T_563 ? 8'h45 : _GEN_4457; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4459 = 8'h69 == _T_563 ? 8'hf9 : _GEN_4458; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4460 = 8'h6a == _T_563 ? 8'h2 : _GEN_4459; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4461 = 8'h6b == _T_563 ? 8'h7f : _GEN_4460; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4462 = 8'h6c == _T_563 ? 8'h50 : _GEN_4461; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4463 = 8'h6d == _T_563 ? 8'h3c : _GEN_4462; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4464 = 8'h6e == _T_563 ? 8'h9f : _GEN_4463; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4465 = 8'h6f == _T_563 ? 8'ha8 : _GEN_4464; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4466 = 8'h70 == _T_563 ? 8'h51 : _GEN_4465; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4467 = 8'h71 == _T_563 ? 8'ha3 : _GEN_4466; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4468 = 8'h72 == _T_563 ? 8'h40 : _GEN_4467; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4469 = 8'h73 == _T_563 ? 8'h8f : _GEN_4468; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4470 = 8'h74 == _T_563 ? 8'h92 : _GEN_4469; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4471 = 8'h75 == _T_563 ? 8'h9d : _GEN_4470; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4472 = 8'h76 == _T_563 ? 8'h38 : _GEN_4471; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4473 = 8'h77 == _T_563 ? 8'hf5 : _GEN_4472; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4474 = 8'h78 == _T_563 ? 8'hbc : _GEN_4473; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4475 = 8'h79 == _T_563 ? 8'hb6 : _GEN_4474; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4476 = 8'h7a == _T_563 ? 8'hda : _GEN_4475; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4477 = 8'h7b == _T_563 ? 8'h21 : _GEN_4476; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4478 = 8'h7c == _T_563 ? 8'h10 : _GEN_4477; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4479 = 8'h7d == _T_563 ? 8'hff : _GEN_4478; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4480 = 8'h7e == _T_563 ? 8'hf3 : _GEN_4479; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4481 = 8'h7f == _T_563 ? 8'hd2 : _GEN_4480; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4482 = 8'h80 == _T_563 ? 8'hcd : _GEN_4481; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4483 = 8'h81 == _T_563 ? 8'hc : _GEN_4482; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4484 = 8'h82 == _T_563 ? 8'h13 : _GEN_4483; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4485 = 8'h83 == _T_563 ? 8'hec : _GEN_4484; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4486 = 8'h84 == _T_563 ? 8'h5f : _GEN_4485; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4487 = 8'h85 == _T_563 ? 8'h97 : _GEN_4486; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4488 = 8'h86 == _T_563 ? 8'h44 : _GEN_4487; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4489 = 8'h87 == _T_563 ? 8'h17 : _GEN_4488; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4490 = 8'h88 == _T_563 ? 8'hc4 : _GEN_4489; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4491 = 8'h89 == _T_563 ? 8'ha7 : _GEN_4490; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4492 = 8'h8a == _T_563 ? 8'h7e : _GEN_4491; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4493 = 8'h8b == _T_563 ? 8'h3d : _GEN_4492; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4494 = 8'h8c == _T_563 ? 8'h64 : _GEN_4493; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4495 = 8'h8d == _T_563 ? 8'h5d : _GEN_4494; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4496 = 8'h8e == _T_563 ? 8'h19 : _GEN_4495; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4497 = 8'h8f == _T_563 ? 8'h73 : _GEN_4496; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4498 = 8'h90 == _T_563 ? 8'h60 : _GEN_4497; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4499 = 8'h91 == _T_563 ? 8'h81 : _GEN_4498; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4500 = 8'h92 == _T_563 ? 8'h4f : _GEN_4499; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4501 = 8'h93 == _T_563 ? 8'hdc : _GEN_4500; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4502 = 8'h94 == _T_563 ? 8'h22 : _GEN_4501; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4503 = 8'h95 == _T_563 ? 8'h2a : _GEN_4502; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4504 = 8'h96 == _T_563 ? 8'h90 : _GEN_4503; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4505 = 8'h97 == _T_563 ? 8'h88 : _GEN_4504; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4506 = 8'h98 == _T_563 ? 8'h46 : _GEN_4505; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4507 = 8'h99 == _T_563 ? 8'hee : _GEN_4506; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4508 = 8'h9a == _T_563 ? 8'hb8 : _GEN_4507; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4509 = 8'h9b == _T_563 ? 8'h14 : _GEN_4508; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4510 = 8'h9c == _T_563 ? 8'hde : _GEN_4509; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4511 = 8'h9d == _T_563 ? 8'h5e : _GEN_4510; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4512 = 8'h9e == _T_563 ? 8'hb : _GEN_4511; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4513 = 8'h9f == _T_563 ? 8'hdb : _GEN_4512; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4514 = 8'ha0 == _T_563 ? 8'he0 : _GEN_4513; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4515 = 8'ha1 == _T_563 ? 8'h32 : _GEN_4514; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4516 = 8'ha2 == _T_563 ? 8'h3a : _GEN_4515; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4517 = 8'ha3 == _T_563 ? 8'ha : _GEN_4516; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4518 = 8'ha4 == _T_563 ? 8'h49 : _GEN_4517; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4519 = 8'ha5 == _T_563 ? 8'h6 : _GEN_4518; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4520 = 8'ha6 == _T_563 ? 8'h24 : _GEN_4519; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4521 = 8'ha7 == _T_563 ? 8'h5c : _GEN_4520; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4522 = 8'ha8 == _T_563 ? 8'hc2 : _GEN_4521; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4523 = 8'ha9 == _T_563 ? 8'hd3 : _GEN_4522; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4524 = 8'haa == _T_563 ? 8'hac : _GEN_4523; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4525 = 8'hab == _T_563 ? 8'h62 : _GEN_4524; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4526 = 8'hac == _T_563 ? 8'h91 : _GEN_4525; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4527 = 8'had == _T_563 ? 8'h95 : _GEN_4526; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4528 = 8'hae == _T_563 ? 8'he4 : _GEN_4527; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4529 = 8'haf == _T_563 ? 8'h79 : _GEN_4528; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4530 = 8'hb0 == _T_563 ? 8'he7 : _GEN_4529; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4531 = 8'hb1 == _T_563 ? 8'hc8 : _GEN_4530; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4532 = 8'hb2 == _T_563 ? 8'h37 : _GEN_4531; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4533 = 8'hb3 == _T_563 ? 8'h6d : _GEN_4532; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4534 = 8'hb4 == _T_563 ? 8'h8d : _GEN_4533; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4535 = 8'hb5 == _T_563 ? 8'hd5 : _GEN_4534; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4536 = 8'hb6 == _T_563 ? 8'h4e : _GEN_4535; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4537 = 8'hb7 == _T_563 ? 8'ha9 : _GEN_4536; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4538 = 8'hb8 == _T_563 ? 8'h6c : _GEN_4537; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4539 = 8'hb9 == _T_563 ? 8'h56 : _GEN_4538; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4540 = 8'hba == _T_563 ? 8'hf4 : _GEN_4539; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4541 = 8'hbb == _T_563 ? 8'hea : _GEN_4540; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4542 = 8'hbc == _T_563 ? 8'h65 : _GEN_4541; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4543 = 8'hbd == _T_563 ? 8'h7a : _GEN_4542; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4544 = 8'hbe == _T_563 ? 8'hae : _GEN_4543; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4545 = 8'hbf == _T_563 ? 8'h8 : _GEN_4544; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4546 = 8'hc0 == _T_563 ? 8'hba : _GEN_4545; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4547 = 8'hc1 == _T_563 ? 8'h78 : _GEN_4546; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4548 = 8'hc2 == _T_563 ? 8'h25 : _GEN_4547; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4549 = 8'hc3 == _T_563 ? 8'h2e : _GEN_4548; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4550 = 8'hc4 == _T_563 ? 8'h1c : _GEN_4549; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4551 = 8'hc5 == _T_563 ? 8'ha6 : _GEN_4550; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4552 = 8'hc6 == _T_563 ? 8'hb4 : _GEN_4551; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4553 = 8'hc7 == _T_563 ? 8'hc6 : _GEN_4552; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4554 = 8'hc8 == _T_563 ? 8'he8 : _GEN_4553; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4555 = 8'hc9 == _T_563 ? 8'hdd : _GEN_4554; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4556 = 8'hca == _T_563 ? 8'h74 : _GEN_4555; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4557 = 8'hcb == _T_563 ? 8'h1f : _GEN_4556; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4558 = 8'hcc == _T_563 ? 8'h4b : _GEN_4557; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4559 = 8'hcd == _T_563 ? 8'hbd : _GEN_4558; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4560 = 8'hce == _T_563 ? 8'h8b : _GEN_4559; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4561 = 8'hcf == _T_563 ? 8'h8a : _GEN_4560; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4562 = 8'hd0 == _T_563 ? 8'h70 : _GEN_4561; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4563 = 8'hd1 == _T_563 ? 8'h3e : _GEN_4562; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4564 = 8'hd2 == _T_563 ? 8'hb5 : _GEN_4563; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4565 = 8'hd3 == _T_563 ? 8'h66 : _GEN_4564; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4566 = 8'hd4 == _T_563 ? 8'h48 : _GEN_4565; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4567 = 8'hd5 == _T_563 ? 8'h3 : _GEN_4566; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4568 = 8'hd6 == _T_563 ? 8'hf6 : _GEN_4567; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4569 = 8'hd7 == _T_563 ? 8'he : _GEN_4568; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4570 = 8'hd8 == _T_563 ? 8'h61 : _GEN_4569; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4571 = 8'hd9 == _T_563 ? 8'h35 : _GEN_4570; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4572 = 8'hda == _T_563 ? 8'h57 : _GEN_4571; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4573 = 8'hdb == _T_563 ? 8'hb9 : _GEN_4572; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4574 = 8'hdc == _T_563 ? 8'h86 : _GEN_4573; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4575 = 8'hdd == _T_563 ? 8'hc1 : _GEN_4574; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4576 = 8'hde == _T_563 ? 8'h1d : _GEN_4575; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4577 = 8'hdf == _T_563 ? 8'h9e : _GEN_4576; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4578 = 8'he0 == _T_563 ? 8'he1 : _GEN_4577; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4579 = 8'he1 == _T_563 ? 8'hf8 : _GEN_4578; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4580 = 8'he2 == _T_563 ? 8'h98 : _GEN_4579; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4581 = 8'he3 == _T_563 ? 8'h11 : _GEN_4580; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4582 = 8'he4 == _T_563 ? 8'h69 : _GEN_4581; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4583 = 8'he5 == _T_563 ? 8'hd9 : _GEN_4582; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4584 = 8'he6 == _T_563 ? 8'h8e : _GEN_4583; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4585 = 8'he7 == _T_563 ? 8'h94 : _GEN_4584; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4586 = 8'he8 == _T_563 ? 8'h9b : _GEN_4585; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4587 = 8'he9 == _T_563 ? 8'h1e : _GEN_4586; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4588 = 8'hea == _T_563 ? 8'h87 : _GEN_4587; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4589 = 8'heb == _T_563 ? 8'he9 : _GEN_4588; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4590 = 8'hec == _T_563 ? 8'hce : _GEN_4589; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4591 = 8'hed == _T_563 ? 8'h55 : _GEN_4590; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4592 = 8'hee == _T_563 ? 8'h28 : _GEN_4591; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4593 = 8'hef == _T_563 ? 8'hdf : _GEN_4592; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4594 = 8'hf0 == _T_563 ? 8'h8c : _GEN_4593; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4595 = 8'hf1 == _T_563 ? 8'ha1 : _GEN_4594; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4596 = 8'hf2 == _T_563 ? 8'h89 : _GEN_4595; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4597 = 8'hf3 == _T_563 ? 8'hd : _GEN_4596; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4598 = 8'hf4 == _T_563 ? 8'hbf : _GEN_4597; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4599 = 8'hf5 == _T_563 ? 8'he6 : _GEN_4598; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4600 = 8'hf6 == _T_563 ? 8'h42 : _GEN_4599; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4601 = 8'hf7 == _T_563 ? 8'h68 : _GEN_4600; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4602 = 8'hf8 == _T_563 ? 8'h41 : _GEN_4601; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4603 = 8'hf9 == _T_563 ? 8'h99 : _GEN_4602; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4604 = 8'hfa == _T_563 ? 8'h2d : _GEN_4603; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4605 = 8'hfb == _T_563 ? 8'hf : _GEN_4604; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4606 = 8'hfc == _T_563 ? 8'hb0 : _GEN_4605; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4607 = 8'hfd == _T_563 ? 8'h54 : _GEN_4606; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4608 = 8'hfe == _T_563 ? 8'hbb : _GEN_4607; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4609 = 8'hff == _T_563 ? 8'h16 : _GEN_4608; // @[Cat.scala 30:58:@2094.4]
  assign _T_571 = {_GEN_4354,_GEN_4609}; // @[Cat.scala 30:58:@2094.4]
  assign _GEN_4610 = 8'h1 == _T_569 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4611 = 8'h2 == _T_569 ? 8'h77 : _GEN_4610; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4612 = 8'h3 == _T_569 ? 8'h7b : _GEN_4611; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4613 = 8'h4 == _T_569 ? 8'hf2 : _GEN_4612; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4614 = 8'h5 == _T_569 ? 8'h6b : _GEN_4613; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4615 = 8'h6 == _T_569 ? 8'h6f : _GEN_4614; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4616 = 8'h7 == _T_569 ? 8'hc5 : _GEN_4615; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4617 = 8'h8 == _T_569 ? 8'h30 : _GEN_4616; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4618 = 8'h9 == _T_569 ? 8'h1 : _GEN_4617; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4619 = 8'ha == _T_569 ? 8'h67 : _GEN_4618; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4620 = 8'hb == _T_569 ? 8'h2b : _GEN_4619; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4621 = 8'hc == _T_569 ? 8'hfe : _GEN_4620; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4622 = 8'hd == _T_569 ? 8'hd7 : _GEN_4621; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4623 = 8'he == _T_569 ? 8'hab : _GEN_4622; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4624 = 8'hf == _T_569 ? 8'h76 : _GEN_4623; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4625 = 8'h10 == _T_569 ? 8'hca : _GEN_4624; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4626 = 8'h11 == _T_569 ? 8'h82 : _GEN_4625; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4627 = 8'h12 == _T_569 ? 8'hc9 : _GEN_4626; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4628 = 8'h13 == _T_569 ? 8'h7d : _GEN_4627; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4629 = 8'h14 == _T_569 ? 8'hfa : _GEN_4628; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4630 = 8'h15 == _T_569 ? 8'h59 : _GEN_4629; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4631 = 8'h16 == _T_569 ? 8'h47 : _GEN_4630; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4632 = 8'h17 == _T_569 ? 8'hf0 : _GEN_4631; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4633 = 8'h18 == _T_569 ? 8'had : _GEN_4632; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4634 = 8'h19 == _T_569 ? 8'hd4 : _GEN_4633; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4635 = 8'h1a == _T_569 ? 8'ha2 : _GEN_4634; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4636 = 8'h1b == _T_569 ? 8'haf : _GEN_4635; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4637 = 8'h1c == _T_569 ? 8'h9c : _GEN_4636; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4638 = 8'h1d == _T_569 ? 8'ha4 : _GEN_4637; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4639 = 8'h1e == _T_569 ? 8'h72 : _GEN_4638; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4640 = 8'h1f == _T_569 ? 8'hc0 : _GEN_4639; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4641 = 8'h20 == _T_569 ? 8'hb7 : _GEN_4640; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4642 = 8'h21 == _T_569 ? 8'hfd : _GEN_4641; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4643 = 8'h22 == _T_569 ? 8'h93 : _GEN_4642; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4644 = 8'h23 == _T_569 ? 8'h26 : _GEN_4643; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4645 = 8'h24 == _T_569 ? 8'h36 : _GEN_4644; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4646 = 8'h25 == _T_569 ? 8'h3f : _GEN_4645; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4647 = 8'h26 == _T_569 ? 8'hf7 : _GEN_4646; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4648 = 8'h27 == _T_569 ? 8'hcc : _GEN_4647; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4649 = 8'h28 == _T_569 ? 8'h34 : _GEN_4648; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4650 = 8'h29 == _T_569 ? 8'ha5 : _GEN_4649; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4651 = 8'h2a == _T_569 ? 8'he5 : _GEN_4650; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4652 = 8'h2b == _T_569 ? 8'hf1 : _GEN_4651; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4653 = 8'h2c == _T_569 ? 8'h71 : _GEN_4652; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4654 = 8'h2d == _T_569 ? 8'hd8 : _GEN_4653; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4655 = 8'h2e == _T_569 ? 8'h31 : _GEN_4654; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4656 = 8'h2f == _T_569 ? 8'h15 : _GEN_4655; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4657 = 8'h30 == _T_569 ? 8'h4 : _GEN_4656; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4658 = 8'h31 == _T_569 ? 8'hc7 : _GEN_4657; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4659 = 8'h32 == _T_569 ? 8'h23 : _GEN_4658; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4660 = 8'h33 == _T_569 ? 8'hc3 : _GEN_4659; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4661 = 8'h34 == _T_569 ? 8'h18 : _GEN_4660; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4662 = 8'h35 == _T_569 ? 8'h96 : _GEN_4661; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4663 = 8'h36 == _T_569 ? 8'h5 : _GEN_4662; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4664 = 8'h37 == _T_569 ? 8'h9a : _GEN_4663; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4665 = 8'h38 == _T_569 ? 8'h7 : _GEN_4664; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4666 = 8'h39 == _T_569 ? 8'h12 : _GEN_4665; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4667 = 8'h3a == _T_569 ? 8'h80 : _GEN_4666; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4668 = 8'h3b == _T_569 ? 8'he2 : _GEN_4667; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4669 = 8'h3c == _T_569 ? 8'heb : _GEN_4668; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4670 = 8'h3d == _T_569 ? 8'h27 : _GEN_4669; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4671 = 8'h3e == _T_569 ? 8'hb2 : _GEN_4670; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4672 = 8'h3f == _T_569 ? 8'h75 : _GEN_4671; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4673 = 8'h40 == _T_569 ? 8'h9 : _GEN_4672; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4674 = 8'h41 == _T_569 ? 8'h83 : _GEN_4673; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4675 = 8'h42 == _T_569 ? 8'h2c : _GEN_4674; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4676 = 8'h43 == _T_569 ? 8'h1a : _GEN_4675; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4677 = 8'h44 == _T_569 ? 8'h1b : _GEN_4676; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4678 = 8'h45 == _T_569 ? 8'h6e : _GEN_4677; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4679 = 8'h46 == _T_569 ? 8'h5a : _GEN_4678; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4680 = 8'h47 == _T_569 ? 8'ha0 : _GEN_4679; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4681 = 8'h48 == _T_569 ? 8'h52 : _GEN_4680; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4682 = 8'h49 == _T_569 ? 8'h3b : _GEN_4681; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4683 = 8'h4a == _T_569 ? 8'hd6 : _GEN_4682; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4684 = 8'h4b == _T_569 ? 8'hb3 : _GEN_4683; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4685 = 8'h4c == _T_569 ? 8'h29 : _GEN_4684; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4686 = 8'h4d == _T_569 ? 8'he3 : _GEN_4685; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4687 = 8'h4e == _T_569 ? 8'h2f : _GEN_4686; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4688 = 8'h4f == _T_569 ? 8'h84 : _GEN_4687; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4689 = 8'h50 == _T_569 ? 8'h53 : _GEN_4688; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4690 = 8'h51 == _T_569 ? 8'hd1 : _GEN_4689; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4691 = 8'h52 == _T_569 ? 8'h0 : _GEN_4690; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4692 = 8'h53 == _T_569 ? 8'hed : _GEN_4691; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4693 = 8'h54 == _T_569 ? 8'h20 : _GEN_4692; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4694 = 8'h55 == _T_569 ? 8'hfc : _GEN_4693; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4695 = 8'h56 == _T_569 ? 8'hb1 : _GEN_4694; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4696 = 8'h57 == _T_569 ? 8'h5b : _GEN_4695; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4697 = 8'h58 == _T_569 ? 8'h6a : _GEN_4696; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4698 = 8'h59 == _T_569 ? 8'hcb : _GEN_4697; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4699 = 8'h5a == _T_569 ? 8'hbe : _GEN_4698; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4700 = 8'h5b == _T_569 ? 8'h39 : _GEN_4699; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4701 = 8'h5c == _T_569 ? 8'h4a : _GEN_4700; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4702 = 8'h5d == _T_569 ? 8'h4c : _GEN_4701; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4703 = 8'h5e == _T_569 ? 8'h58 : _GEN_4702; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4704 = 8'h5f == _T_569 ? 8'hcf : _GEN_4703; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4705 = 8'h60 == _T_569 ? 8'hd0 : _GEN_4704; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4706 = 8'h61 == _T_569 ? 8'hef : _GEN_4705; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4707 = 8'h62 == _T_569 ? 8'haa : _GEN_4706; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4708 = 8'h63 == _T_569 ? 8'hfb : _GEN_4707; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4709 = 8'h64 == _T_569 ? 8'h43 : _GEN_4708; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4710 = 8'h65 == _T_569 ? 8'h4d : _GEN_4709; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4711 = 8'h66 == _T_569 ? 8'h33 : _GEN_4710; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4712 = 8'h67 == _T_569 ? 8'h85 : _GEN_4711; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4713 = 8'h68 == _T_569 ? 8'h45 : _GEN_4712; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4714 = 8'h69 == _T_569 ? 8'hf9 : _GEN_4713; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4715 = 8'h6a == _T_569 ? 8'h2 : _GEN_4714; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4716 = 8'h6b == _T_569 ? 8'h7f : _GEN_4715; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4717 = 8'h6c == _T_569 ? 8'h50 : _GEN_4716; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4718 = 8'h6d == _T_569 ? 8'h3c : _GEN_4717; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4719 = 8'h6e == _T_569 ? 8'h9f : _GEN_4718; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4720 = 8'h6f == _T_569 ? 8'ha8 : _GEN_4719; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4721 = 8'h70 == _T_569 ? 8'h51 : _GEN_4720; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4722 = 8'h71 == _T_569 ? 8'ha3 : _GEN_4721; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4723 = 8'h72 == _T_569 ? 8'h40 : _GEN_4722; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4724 = 8'h73 == _T_569 ? 8'h8f : _GEN_4723; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4725 = 8'h74 == _T_569 ? 8'h92 : _GEN_4724; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4726 = 8'h75 == _T_569 ? 8'h9d : _GEN_4725; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4727 = 8'h76 == _T_569 ? 8'h38 : _GEN_4726; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4728 = 8'h77 == _T_569 ? 8'hf5 : _GEN_4727; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4729 = 8'h78 == _T_569 ? 8'hbc : _GEN_4728; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4730 = 8'h79 == _T_569 ? 8'hb6 : _GEN_4729; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4731 = 8'h7a == _T_569 ? 8'hda : _GEN_4730; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4732 = 8'h7b == _T_569 ? 8'h21 : _GEN_4731; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4733 = 8'h7c == _T_569 ? 8'h10 : _GEN_4732; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4734 = 8'h7d == _T_569 ? 8'hff : _GEN_4733; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4735 = 8'h7e == _T_569 ? 8'hf3 : _GEN_4734; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4736 = 8'h7f == _T_569 ? 8'hd2 : _GEN_4735; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4737 = 8'h80 == _T_569 ? 8'hcd : _GEN_4736; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4738 = 8'h81 == _T_569 ? 8'hc : _GEN_4737; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4739 = 8'h82 == _T_569 ? 8'h13 : _GEN_4738; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4740 = 8'h83 == _T_569 ? 8'hec : _GEN_4739; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4741 = 8'h84 == _T_569 ? 8'h5f : _GEN_4740; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4742 = 8'h85 == _T_569 ? 8'h97 : _GEN_4741; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4743 = 8'h86 == _T_569 ? 8'h44 : _GEN_4742; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4744 = 8'h87 == _T_569 ? 8'h17 : _GEN_4743; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4745 = 8'h88 == _T_569 ? 8'hc4 : _GEN_4744; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4746 = 8'h89 == _T_569 ? 8'ha7 : _GEN_4745; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4747 = 8'h8a == _T_569 ? 8'h7e : _GEN_4746; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4748 = 8'h8b == _T_569 ? 8'h3d : _GEN_4747; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4749 = 8'h8c == _T_569 ? 8'h64 : _GEN_4748; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4750 = 8'h8d == _T_569 ? 8'h5d : _GEN_4749; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4751 = 8'h8e == _T_569 ? 8'h19 : _GEN_4750; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4752 = 8'h8f == _T_569 ? 8'h73 : _GEN_4751; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4753 = 8'h90 == _T_569 ? 8'h60 : _GEN_4752; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4754 = 8'h91 == _T_569 ? 8'h81 : _GEN_4753; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4755 = 8'h92 == _T_569 ? 8'h4f : _GEN_4754; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4756 = 8'h93 == _T_569 ? 8'hdc : _GEN_4755; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4757 = 8'h94 == _T_569 ? 8'h22 : _GEN_4756; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4758 = 8'h95 == _T_569 ? 8'h2a : _GEN_4757; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4759 = 8'h96 == _T_569 ? 8'h90 : _GEN_4758; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4760 = 8'h97 == _T_569 ? 8'h88 : _GEN_4759; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4761 = 8'h98 == _T_569 ? 8'h46 : _GEN_4760; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4762 = 8'h99 == _T_569 ? 8'hee : _GEN_4761; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4763 = 8'h9a == _T_569 ? 8'hb8 : _GEN_4762; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4764 = 8'h9b == _T_569 ? 8'h14 : _GEN_4763; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4765 = 8'h9c == _T_569 ? 8'hde : _GEN_4764; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4766 = 8'h9d == _T_569 ? 8'h5e : _GEN_4765; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4767 = 8'h9e == _T_569 ? 8'hb : _GEN_4766; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4768 = 8'h9f == _T_569 ? 8'hdb : _GEN_4767; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4769 = 8'ha0 == _T_569 ? 8'he0 : _GEN_4768; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4770 = 8'ha1 == _T_569 ? 8'h32 : _GEN_4769; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4771 = 8'ha2 == _T_569 ? 8'h3a : _GEN_4770; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4772 = 8'ha3 == _T_569 ? 8'ha : _GEN_4771; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4773 = 8'ha4 == _T_569 ? 8'h49 : _GEN_4772; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4774 = 8'ha5 == _T_569 ? 8'h6 : _GEN_4773; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4775 = 8'ha6 == _T_569 ? 8'h24 : _GEN_4774; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4776 = 8'ha7 == _T_569 ? 8'h5c : _GEN_4775; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4777 = 8'ha8 == _T_569 ? 8'hc2 : _GEN_4776; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4778 = 8'ha9 == _T_569 ? 8'hd3 : _GEN_4777; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4779 = 8'haa == _T_569 ? 8'hac : _GEN_4778; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4780 = 8'hab == _T_569 ? 8'h62 : _GEN_4779; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4781 = 8'hac == _T_569 ? 8'h91 : _GEN_4780; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4782 = 8'had == _T_569 ? 8'h95 : _GEN_4781; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4783 = 8'hae == _T_569 ? 8'he4 : _GEN_4782; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4784 = 8'haf == _T_569 ? 8'h79 : _GEN_4783; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4785 = 8'hb0 == _T_569 ? 8'he7 : _GEN_4784; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4786 = 8'hb1 == _T_569 ? 8'hc8 : _GEN_4785; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4787 = 8'hb2 == _T_569 ? 8'h37 : _GEN_4786; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4788 = 8'hb3 == _T_569 ? 8'h6d : _GEN_4787; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4789 = 8'hb4 == _T_569 ? 8'h8d : _GEN_4788; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4790 = 8'hb5 == _T_569 ? 8'hd5 : _GEN_4789; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4791 = 8'hb6 == _T_569 ? 8'h4e : _GEN_4790; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4792 = 8'hb7 == _T_569 ? 8'ha9 : _GEN_4791; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4793 = 8'hb8 == _T_569 ? 8'h6c : _GEN_4792; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4794 = 8'hb9 == _T_569 ? 8'h56 : _GEN_4793; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4795 = 8'hba == _T_569 ? 8'hf4 : _GEN_4794; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4796 = 8'hbb == _T_569 ? 8'hea : _GEN_4795; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4797 = 8'hbc == _T_569 ? 8'h65 : _GEN_4796; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4798 = 8'hbd == _T_569 ? 8'h7a : _GEN_4797; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4799 = 8'hbe == _T_569 ? 8'hae : _GEN_4798; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4800 = 8'hbf == _T_569 ? 8'h8 : _GEN_4799; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4801 = 8'hc0 == _T_569 ? 8'hba : _GEN_4800; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4802 = 8'hc1 == _T_569 ? 8'h78 : _GEN_4801; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4803 = 8'hc2 == _T_569 ? 8'h25 : _GEN_4802; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4804 = 8'hc3 == _T_569 ? 8'h2e : _GEN_4803; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4805 = 8'hc4 == _T_569 ? 8'h1c : _GEN_4804; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4806 = 8'hc5 == _T_569 ? 8'ha6 : _GEN_4805; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4807 = 8'hc6 == _T_569 ? 8'hb4 : _GEN_4806; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4808 = 8'hc7 == _T_569 ? 8'hc6 : _GEN_4807; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4809 = 8'hc8 == _T_569 ? 8'he8 : _GEN_4808; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4810 = 8'hc9 == _T_569 ? 8'hdd : _GEN_4809; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4811 = 8'hca == _T_569 ? 8'h74 : _GEN_4810; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4812 = 8'hcb == _T_569 ? 8'h1f : _GEN_4811; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4813 = 8'hcc == _T_569 ? 8'h4b : _GEN_4812; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4814 = 8'hcd == _T_569 ? 8'hbd : _GEN_4813; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4815 = 8'hce == _T_569 ? 8'h8b : _GEN_4814; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4816 = 8'hcf == _T_569 ? 8'h8a : _GEN_4815; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4817 = 8'hd0 == _T_569 ? 8'h70 : _GEN_4816; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4818 = 8'hd1 == _T_569 ? 8'h3e : _GEN_4817; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4819 = 8'hd2 == _T_569 ? 8'hb5 : _GEN_4818; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4820 = 8'hd3 == _T_569 ? 8'h66 : _GEN_4819; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4821 = 8'hd4 == _T_569 ? 8'h48 : _GEN_4820; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4822 = 8'hd5 == _T_569 ? 8'h3 : _GEN_4821; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4823 = 8'hd6 == _T_569 ? 8'hf6 : _GEN_4822; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4824 = 8'hd7 == _T_569 ? 8'he : _GEN_4823; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4825 = 8'hd8 == _T_569 ? 8'h61 : _GEN_4824; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4826 = 8'hd9 == _T_569 ? 8'h35 : _GEN_4825; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4827 = 8'hda == _T_569 ? 8'h57 : _GEN_4826; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4828 = 8'hdb == _T_569 ? 8'hb9 : _GEN_4827; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4829 = 8'hdc == _T_569 ? 8'h86 : _GEN_4828; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4830 = 8'hdd == _T_569 ? 8'hc1 : _GEN_4829; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4831 = 8'hde == _T_569 ? 8'h1d : _GEN_4830; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4832 = 8'hdf == _T_569 ? 8'h9e : _GEN_4831; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4833 = 8'he0 == _T_569 ? 8'he1 : _GEN_4832; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4834 = 8'he1 == _T_569 ? 8'hf8 : _GEN_4833; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4835 = 8'he2 == _T_569 ? 8'h98 : _GEN_4834; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4836 = 8'he3 == _T_569 ? 8'h11 : _GEN_4835; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4837 = 8'he4 == _T_569 ? 8'h69 : _GEN_4836; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4838 = 8'he5 == _T_569 ? 8'hd9 : _GEN_4837; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4839 = 8'he6 == _T_569 ? 8'h8e : _GEN_4838; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4840 = 8'he7 == _T_569 ? 8'h94 : _GEN_4839; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4841 = 8'he8 == _T_569 ? 8'h9b : _GEN_4840; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4842 = 8'he9 == _T_569 ? 8'h1e : _GEN_4841; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4843 = 8'hea == _T_569 ? 8'h87 : _GEN_4842; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4844 = 8'heb == _T_569 ? 8'he9 : _GEN_4843; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4845 = 8'hec == _T_569 ? 8'hce : _GEN_4844; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4846 = 8'hed == _T_569 ? 8'h55 : _GEN_4845; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4847 = 8'hee == _T_569 ? 8'h28 : _GEN_4846; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4848 = 8'hef == _T_569 ? 8'hdf : _GEN_4847; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4849 = 8'hf0 == _T_569 ? 8'h8c : _GEN_4848; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4850 = 8'hf1 == _T_569 ? 8'ha1 : _GEN_4849; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4851 = 8'hf2 == _T_569 ? 8'h89 : _GEN_4850; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4852 = 8'hf3 == _T_569 ? 8'hd : _GEN_4851; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4853 = 8'hf4 == _T_569 ? 8'hbf : _GEN_4852; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4854 = 8'hf5 == _T_569 ? 8'he6 : _GEN_4853; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4855 = 8'hf6 == _T_569 ? 8'h42 : _GEN_4854; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4856 = 8'hf7 == _T_569 ? 8'h68 : _GEN_4855; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4857 = 8'hf8 == _T_569 ? 8'h41 : _GEN_4856; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4858 = 8'hf9 == _T_569 ? 8'h99 : _GEN_4857; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4859 = 8'hfa == _T_569 ? 8'h2d : _GEN_4858; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4860 = 8'hfb == _T_569 ? 8'hf : _GEN_4859; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4861 = 8'hfc == _T_569 ? 8'hb0 : _GEN_4860; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4862 = 8'hfd == _T_569 ? 8'h54 : _GEN_4861; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4863 = 8'hfe == _T_569 ? 8'hbb : _GEN_4862; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4864 = 8'hff == _T_569 ? 8'h16 : _GEN_4863; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4865 = 8'h1 == _T_567 ? 8'h7c : 8'h63; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4866 = 8'h2 == _T_567 ? 8'h77 : _GEN_4865; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4867 = 8'h3 == _T_567 ? 8'h7b : _GEN_4866; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4868 = 8'h4 == _T_567 ? 8'hf2 : _GEN_4867; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4869 = 8'h5 == _T_567 ? 8'h6b : _GEN_4868; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4870 = 8'h6 == _T_567 ? 8'h6f : _GEN_4869; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4871 = 8'h7 == _T_567 ? 8'hc5 : _GEN_4870; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4872 = 8'h8 == _T_567 ? 8'h30 : _GEN_4871; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4873 = 8'h9 == _T_567 ? 8'h1 : _GEN_4872; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4874 = 8'ha == _T_567 ? 8'h67 : _GEN_4873; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4875 = 8'hb == _T_567 ? 8'h2b : _GEN_4874; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4876 = 8'hc == _T_567 ? 8'hfe : _GEN_4875; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4877 = 8'hd == _T_567 ? 8'hd7 : _GEN_4876; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4878 = 8'he == _T_567 ? 8'hab : _GEN_4877; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4879 = 8'hf == _T_567 ? 8'h76 : _GEN_4878; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4880 = 8'h10 == _T_567 ? 8'hca : _GEN_4879; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4881 = 8'h11 == _T_567 ? 8'h82 : _GEN_4880; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4882 = 8'h12 == _T_567 ? 8'hc9 : _GEN_4881; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4883 = 8'h13 == _T_567 ? 8'h7d : _GEN_4882; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4884 = 8'h14 == _T_567 ? 8'hfa : _GEN_4883; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4885 = 8'h15 == _T_567 ? 8'h59 : _GEN_4884; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4886 = 8'h16 == _T_567 ? 8'h47 : _GEN_4885; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4887 = 8'h17 == _T_567 ? 8'hf0 : _GEN_4886; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4888 = 8'h18 == _T_567 ? 8'had : _GEN_4887; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4889 = 8'h19 == _T_567 ? 8'hd4 : _GEN_4888; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4890 = 8'h1a == _T_567 ? 8'ha2 : _GEN_4889; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4891 = 8'h1b == _T_567 ? 8'haf : _GEN_4890; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4892 = 8'h1c == _T_567 ? 8'h9c : _GEN_4891; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4893 = 8'h1d == _T_567 ? 8'ha4 : _GEN_4892; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4894 = 8'h1e == _T_567 ? 8'h72 : _GEN_4893; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4895 = 8'h1f == _T_567 ? 8'hc0 : _GEN_4894; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4896 = 8'h20 == _T_567 ? 8'hb7 : _GEN_4895; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4897 = 8'h21 == _T_567 ? 8'hfd : _GEN_4896; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4898 = 8'h22 == _T_567 ? 8'h93 : _GEN_4897; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4899 = 8'h23 == _T_567 ? 8'h26 : _GEN_4898; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4900 = 8'h24 == _T_567 ? 8'h36 : _GEN_4899; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4901 = 8'h25 == _T_567 ? 8'h3f : _GEN_4900; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4902 = 8'h26 == _T_567 ? 8'hf7 : _GEN_4901; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4903 = 8'h27 == _T_567 ? 8'hcc : _GEN_4902; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4904 = 8'h28 == _T_567 ? 8'h34 : _GEN_4903; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4905 = 8'h29 == _T_567 ? 8'ha5 : _GEN_4904; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4906 = 8'h2a == _T_567 ? 8'he5 : _GEN_4905; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4907 = 8'h2b == _T_567 ? 8'hf1 : _GEN_4906; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4908 = 8'h2c == _T_567 ? 8'h71 : _GEN_4907; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4909 = 8'h2d == _T_567 ? 8'hd8 : _GEN_4908; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4910 = 8'h2e == _T_567 ? 8'h31 : _GEN_4909; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4911 = 8'h2f == _T_567 ? 8'h15 : _GEN_4910; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4912 = 8'h30 == _T_567 ? 8'h4 : _GEN_4911; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4913 = 8'h31 == _T_567 ? 8'hc7 : _GEN_4912; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4914 = 8'h32 == _T_567 ? 8'h23 : _GEN_4913; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4915 = 8'h33 == _T_567 ? 8'hc3 : _GEN_4914; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4916 = 8'h34 == _T_567 ? 8'h18 : _GEN_4915; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4917 = 8'h35 == _T_567 ? 8'h96 : _GEN_4916; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4918 = 8'h36 == _T_567 ? 8'h5 : _GEN_4917; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4919 = 8'h37 == _T_567 ? 8'h9a : _GEN_4918; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4920 = 8'h38 == _T_567 ? 8'h7 : _GEN_4919; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4921 = 8'h39 == _T_567 ? 8'h12 : _GEN_4920; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4922 = 8'h3a == _T_567 ? 8'h80 : _GEN_4921; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4923 = 8'h3b == _T_567 ? 8'he2 : _GEN_4922; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4924 = 8'h3c == _T_567 ? 8'heb : _GEN_4923; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4925 = 8'h3d == _T_567 ? 8'h27 : _GEN_4924; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4926 = 8'h3e == _T_567 ? 8'hb2 : _GEN_4925; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4927 = 8'h3f == _T_567 ? 8'h75 : _GEN_4926; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4928 = 8'h40 == _T_567 ? 8'h9 : _GEN_4927; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4929 = 8'h41 == _T_567 ? 8'h83 : _GEN_4928; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4930 = 8'h42 == _T_567 ? 8'h2c : _GEN_4929; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4931 = 8'h43 == _T_567 ? 8'h1a : _GEN_4930; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4932 = 8'h44 == _T_567 ? 8'h1b : _GEN_4931; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4933 = 8'h45 == _T_567 ? 8'h6e : _GEN_4932; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4934 = 8'h46 == _T_567 ? 8'h5a : _GEN_4933; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4935 = 8'h47 == _T_567 ? 8'ha0 : _GEN_4934; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4936 = 8'h48 == _T_567 ? 8'h52 : _GEN_4935; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4937 = 8'h49 == _T_567 ? 8'h3b : _GEN_4936; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4938 = 8'h4a == _T_567 ? 8'hd6 : _GEN_4937; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4939 = 8'h4b == _T_567 ? 8'hb3 : _GEN_4938; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4940 = 8'h4c == _T_567 ? 8'h29 : _GEN_4939; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4941 = 8'h4d == _T_567 ? 8'he3 : _GEN_4940; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4942 = 8'h4e == _T_567 ? 8'h2f : _GEN_4941; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4943 = 8'h4f == _T_567 ? 8'h84 : _GEN_4942; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4944 = 8'h50 == _T_567 ? 8'h53 : _GEN_4943; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4945 = 8'h51 == _T_567 ? 8'hd1 : _GEN_4944; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4946 = 8'h52 == _T_567 ? 8'h0 : _GEN_4945; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4947 = 8'h53 == _T_567 ? 8'hed : _GEN_4946; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4948 = 8'h54 == _T_567 ? 8'h20 : _GEN_4947; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4949 = 8'h55 == _T_567 ? 8'hfc : _GEN_4948; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4950 = 8'h56 == _T_567 ? 8'hb1 : _GEN_4949; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4951 = 8'h57 == _T_567 ? 8'h5b : _GEN_4950; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4952 = 8'h58 == _T_567 ? 8'h6a : _GEN_4951; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4953 = 8'h59 == _T_567 ? 8'hcb : _GEN_4952; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4954 = 8'h5a == _T_567 ? 8'hbe : _GEN_4953; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4955 = 8'h5b == _T_567 ? 8'h39 : _GEN_4954; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4956 = 8'h5c == _T_567 ? 8'h4a : _GEN_4955; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4957 = 8'h5d == _T_567 ? 8'h4c : _GEN_4956; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4958 = 8'h5e == _T_567 ? 8'h58 : _GEN_4957; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4959 = 8'h5f == _T_567 ? 8'hcf : _GEN_4958; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4960 = 8'h60 == _T_567 ? 8'hd0 : _GEN_4959; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4961 = 8'h61 == _T_567 ? 8'hef : _GEN_4960; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4962 = 8'h62 == _T_567 ? 8'haa : _GEN_4961; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4963 = 8'h63 == _T_567 ? 8'hfb : _GEN_4962; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4964 = 8'h64 == _T_567 ? 8'h43 : _GEN_4963; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4965 = 8'h65 == _T_567 ? 8'h4d : _GEN_4964; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4966 = 8'h66 == _T_567 ? 8'h33 : _GEN_4965; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4967 = 8'h67 == _T_567 ? 8'h85 : _GEN_4966; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4968 = 8'h68 == _T_567 ? 8'h45 : _GEN_4967; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4969 = 8'h69 == _T_567 ? 8'hf9 : _GEN_4968; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4970 = 8'h6a == _T_567 ? 8'h2 : _GEN_4969; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4971 = 8'h6b == _T_567 ? 8'h7f : _GEN_4970; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4972 = 8'h6c == _T_567 ? 8'h50 : _GEN_4971; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4973 = 8'h6d == _T_567 ? 8'h3c : _GEN_4972; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4974 = 8'h6e == _T_567 ? 8'h9f : _GEN_4973; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4975 = 8'h6f == _T_567 ? 8'ha8 : _GEN_4974; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4976 = 8'h70 == _T_567 ? 8'h51 : _GEN_4975; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4977 = 8'h71 == _T_567 ? 8'ha3 : _GEN_4976; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4978 = 8'h72 == _T_567 ? 8'h40 : _GEN_4977; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4979 = 8'h73 == _T_567 ? 8'h8f : _GEN_4978; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4980 = 8'h74 == _T_567 ? 8'h92 : _GEN_4979; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4981 = 8'h75 == _T_567 ? 8'h9d : _GEN_4980; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4982 = 8'h76 == _T_567 ? 8'h38 : _GEN_4981; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4983 = 8'h77 == _T_567 ? 8'hf5 : _GEN_4982; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4984 = 8'h78 == _T_567 ? 8'hbc : _GEN_4983; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4985 = 8'h79 == _T_567 ? 8'hb6 : _GEN_4984; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4986 = 8'h7a == _T_567 ? 8'hda : _GEN_4985; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4987 = 8'h7b == _T_567 ? 8'h21 : _GEN_4986; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4988 = 8'h7c == _T_567 ? 8'h10 : _GEN_4987; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4989 = 8'h7d == _T_567 ? 8'hff : _GEN_4988; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4990 = 8'h7e == _T_567 ? 8'hf3 : _GEN_4989; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4991 = 8'h7f == _T_567 ? 8'hd2 : _GEN_4990; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4992 = 8'h80 == _T_567 ? 8'hcd : _GEN_4991; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4993 = 8'h81 == _T_567 ? 8'hc : _GEN_4992; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4994 = 8'h82 == _T_567 ? 8'h13 : _GEN_4993; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4995 = 8'h83 == _T_567 ? 8'hec : _GEN_4994; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4996 = 8'h84 == _T_567 ? 8'h5f : _GEN_4995; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4997 = 8'h85 == _T_567 ? 8'h97 : _GEN_4996; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4998 = 8'h86 == _T_567 ? 8'h44 : _GEN_4997; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_4999 = 8'h87 == _T_567 ? 8'h17 : _GEN_4998; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5000 = 8'h88 == _T_567 ? 8'hc4 : _GEN_4999; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5001 = 8'h89 == _T_567 ? 8'ha7 : _GEN_5000; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5002 = 8'h8a == _T_567 ? 8'h7e : _GEN_5001; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5003 = 8'h8b == _T_567 ? 8'h3d : _GEN_5002; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5004 = 8'h8c == _T_567 ? 8'h64 : _GEN_5003; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5005 = 8'h8d == _T_567 ? 8'h5d : _GEN_5004; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5006 = 8'h8e == _T_567 ? 8'h19 : _GEN_5005; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5007 = 8'h8f == _T_567 ? 8'h73 : _GEN_5006; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5008 = 8'h90 == _T_567 ? 8'h60 : _GEN_5007; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5009 = 8'h91 == _T_567 ? 8'h81 : _GEN_5008; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5010 = 8'h92 == _T_567 ? 8'h4f : _GEN_5009; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5011 = 8'h93 == _T_567 ? 8'hdc : _GEN_5010; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5012 = 8'h94 == _T_567 ? 8'h22 : _GEN_5011; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5013 = 8'h95 == _T_567 ? 8'h2a : _GEN_5012; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5014 = 8'h96 == _T_567 ? 8'h90 : _GEN_5013; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5015 = 8'h97 == _T_567 ? 8'h88 : _GEN_5014; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5016 = 8'h98 == _T_567 ? 8'h46 : _GEN_5015; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5017 = 8'h99 == _T_567 ? 8'hee : _GEN_5016; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5018 = 8'h9a == _T_567 ? 8'hb8 : _GEN_5017; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5019 = 8'h9b == _T_567 ? 8'h14 : _GEN_5018; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5020 = 8'h9c == _T_567 ? 8'hde : _GEN_5019; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5021 = 8'h9d == _T_567 ? 8'h5e : _GEN_5020; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5022 = 8'h9e == _T_567 ? 8'hb : _GEN_5021; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5023 = 8'h9f == _T_567 ? 8'hdb : _GEN_5022; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5024 = 8'ha0 == _T_567 ? 8'he0 : _GEN_5023; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5025 = 8'ha1 == _T_567 ? 8'h32 : _GEN_5024; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5026 = 8'ha2 == _T_567 ? 8'h3a : _GEN_5025; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5027 = 8'ha3 == _T_567 ? 8'ha : _GEN_5026; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5028 = 8'ha4 == _T_567 ? 8'h49 : _GEN_5027; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5029 = 8'ha5 == _T_567 ? 8'h6 : _GEN_5028; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5030 = 8'ha6 == _T_567 ? 8'h24 : _GEN_5029; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5031 = 8'ha7 == _T_567 ? 8'h5c : _GEN_5030; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5032 = 8'ha8 == _T_567 ? 8'hc2 : _GEN_5031; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5033 = 8'ha9 == _T_567 ? 8'hd3 : _GEN_5032; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5034 = 8'haa == _T_567 ? 8'hac : _GEN_5033; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5035 = 8'hab == _T_567 ? 8'h62 : _GEN_5034; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5036 = 8'hac == _T_567 ? 8'h91 : _GEN_5035; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5037 = 8'had == _T_567 ? 8'h95 : _GEN_5036; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5038 = 8'hae == _T_567 ? 8'he4 : _GEN_5037; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5039 = 8'haf == _T_567 ? 8'h79 : _GEN_5038; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5040 = 8'hb0 == _T_567 ? 8'he7 : _GEN_5039; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5041 = 8'hb1 == _T_567 ? 8'hc8 : _GEN_5040; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5042 = 8'hb2 == _T_567 ? 8'h37 : _GEN_5041; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5043 = 8'hb3 == _T_567 ? 8'h6d : _GEN_5042; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5044 = 8'hb4 == _T_567 ? 8'h8d : _GEN_5043; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5045 = 8'hb5 == _T_567 ? 8'hd5 : _GEN_5044; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5046 = 8'hb6 == _T_567 ? 8'h4e : _GEN_5045; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5047 = 8'hb7 == _T_567 ? 8'ha9 : _GEN_5046; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5048 = 8'hb8 == _T_567 ? 8'h6c : _GEN_5047; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5049 = 8'hb9 == _T_567 ? 8'h56 : _GEN_5048; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5050 = 8'hba == _T_567 ? 8'hf4 : _GEN_5049; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5051 = 8'hbb == _T_567 ? 8'hea : _GEN_5050; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5052 = 8'hbc == _T_567 ? 8'h65 : _GEN_5051; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5053 = 8'hbd == _T_567 ? 8'h7a : _GEN_5052; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5054 = 8'hbe == _T_567 ? 8'hae : _GEN_5053; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5055 = 8'hbf == _T_567 ? 8'h8 : _GEN_5054; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5056 = 8'hc0 == _T_567 ? 8'hba : _GEN_5055; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5057 = 8'hc1 == _T_567 ? 8'h78 : _GEN_5056; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5058 = 8'hc2 == _T_567 ? 8'h25 : _GEN_5057; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5059 = 8'hc3 == _T_567 ? 8'h2e : _GEN_5058; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5060 = 8'hc4 == _T_567 ? 8'h1c : _GEN_5059; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5061 = 8'hc5 == _T_567 ? 8'ha6 : _GEN_5060; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5062 = 8'hc6 == _T_567 ? 8'hb4 : _GEN_5061; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5063 = 8'hc7 == _T_567 ? 8'hc6 : _GEN_5062; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5064 = 8'hc8 == _T_567 ? 8'he8 : _GEN_5063; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5065 = 8'hc9 == _T_567 ? 8'hdd : _GEN_5064; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5066 = 8'hca == _T_567 ? 8'h74 : _GEN_5065; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5067 = 8'hcb == _T_567 ? 8'h1f : _GEN_5066; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5068 = 8'hcc == _T_567 ? 8'h4b : _GEN_5067; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5069 = 8'hcd == _T_567 ? 8'hbd : _GEN_5068; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5070 = 8'hce == _T_567 ? 8'h8b : _GEN_5069; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5071 = 8'hcf == _T_567 ? 8'h8a : _GEN_5070; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5072 = 8'hd0 == _T_567 ? 8'h70 : _GEN_5071; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5073 = 8'hd1 == _T_567 ? 8'h3e : _GEN_5072; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5074 = 8'hd2 == _T_567 ? 8'hb5 : _GEN_5073; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5075 = 8'hd3 == _T_567 ? 8'h66 : _GEN_5074; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5076 = 8'hd4 == _T_567 ? 8'h48 : _GEN_5075; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5077 = 8'hd5 == _T_567 ? 8'h3 : _GEN_5076; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5078 = 8'hd6 == _T_567 ? 8'hf6 : _GEN_5077; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5079 = 8'hd7 == _T_567 ? 8'he : _GEN_5078; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5080 = 8'hd8 == _T_567 ? 8'h61 : _GEN_5079; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5081 = 8'hd9 == _T_567 ? 8'h35 : _GEN_5080; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5082 = 8'hda == _T_567 ? 8'h57 : _GEN_5081; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5083 = 8'hdb == _T_567 ? 8'hb9 : _GEN_5082; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5084 = 8'hdc == _T_567 ? 8'h86 : _GEN_5083; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5085 = 8'hdd == _T_567 ? 8'hc1 : _GEN_5084; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5086 = 8'hde == _T_567 ? 8'h1d : _GEN_5085; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5087 = 8'hdf == _T_567 ? 8'h9e : _GEN_5086; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5088 = 8'he0 == _T_567 ? 8'he1 : _GEN_5087; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5089 = 8'he1 == _T_567 ? 8'hf8 : _GEN_5088; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5090 = 8'he2 == _T_567 ? 8'h98 : _GEN_5089; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5091 = 8'he3 == _T_567 ? 8'h11 : _GEN_5090; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5092 = 8'he4 == _T_567 ? 8'h69 : _GEN_5091; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5093 = 8'he5 == _T_567 ? 8'hd9 : _GEN_5092; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5094 = 8'he6 == _T_567 ? 8'h8e : _GEN_5093; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5095 = 8'he7 == _T_567 ? 8'h94 : _GEN_5094; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5096 = 8'he8 == _T_567 ? 8'h9b : _GEN_5095; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5097 = 8'he9 == _T_567 ? 8'h1e : _GEN_5096; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5098 = 8'hea == _T_567 ? 8'h87 : _GEN_5097; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5099 = 8'heb == _T_567 ? 8'he9 : _GEN_5098; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5100 = 8'hec == _T_567 ? 8'hce : _GEN_5099; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5101 = 8'hed == _T_567 ? 8'h55 : _GEN_5100; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5102 = 8'hee == _T_567 ? 8'h28 : _GEN_5101; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5103 = 8'hef == _T_567 ? 8'hdf : _GEN_5102; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5104 = 8'hf0 == _T_567 ? 8'h8c : _GEN_5103; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5105 = 8'hf1 == _T_567 ? 8'ha1 : _GEN_5104; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5106 = 8'hf2 == _T_567 ? 8'h89 : _GEN_5105; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5107 = 8'hf3 == _T_567 ? 8'hd : _GEN_5106; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5108 = 8'hf4 == _T_567 ? 8'hbf : _GEN_5107; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5109 = 8'hf5 == _T_567 ? 8'he6 : _GEN_5108; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5110 = 8'hf6 == _T_567 ? 8'h42 : _GEN_5109; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5111 = 8'hf7 == _T_567 ? 8'h68 : _GEN_5110; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5112 = 8'hf8 == _T_567 ? 8'h41 : _GEN_5111; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5113 = 8'hf9 == _T_567 ? 8'h99 : _GEN_5112; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5114 = 8'hfa == _T_567 ? 8'h2d : _GEN_5113; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5115 = 8'hfb == _T_567 ? 8'hf : _GEN_5114; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5116 = 8'hfc == _T_567 ? 8'hb0 : _GEN_5115; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5117 = 8'hfd == _T_567 ? 8'h54 : _GEN_5116; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5118 = 8'hfe == _T_567 ? 8'hbb : _GEN_5117; // @[Cat.scala 30:58:@2095.4]
  assign _GEN_5119 = 8'hff == _T_567 ? 8'h16 : _GEN_5118; // @[Cat.scala 30:58:@2095.4]
  assign _T_572 = {_GEN_4864,_GEN_5119}; // @[Cat.scala 30:58:@2095.4]
  assign x4 = {_T_572,_T_571}; // @[Cat.scala 30:58:@2096.4]
  assign _T_573 = {x2,x1}; // @[Cat.scala 30:58:@2097.4]
  assign _T_574 = {x4,x3}; // @[Cat.scala 30:58:@2098.4]
  assign _T_575 = {_T_574,_T_573}; // @[Cat.scala 30:58:@2099.4]
  assign io_data = _T_532;
  assign io_data2 = _T_575;
endmodule
module aes( // @[:@2102.2]
  input          clock, // @[:@2103.4]
  input          reset, // @[:@2104.4]
  output [127:0] io_result, // @[:@2105.4]
  input  [127:0] io_iData, // @[:@2105.4]
  input  [127:0] io_key, // @[:@2105.4]
  output         io_done, // @[:@2105.4]
  input          io_en // @[:@2105.4]
);
  wire  encm_clock; // @[aes.scala 20:19:@2107.4]
  wire  encm_reset; // @[aes.scala 20:19:@2107.4]
  wire [127:0] encm_io_rkey; // @[aes.scala 20:19:@2107.4]
  wire  encm_io_done; // @[aes.scala 20:19:@2107.4]
  wire [127:0] encm_io_sio_addr2; // @[aes.scala 20:19:@2107.4]
  wire [127:0] encm_io_sio_data2; // @[aes.scala 20:19:@2107.4]
  wire [127:0] encm_io_out; // @[aes.scala 20:19:@2107.4]
  wire [3:0] encm_io_roundOut; // @[aes.scala 20:19:@2107.4]
  wire [127:0] encm_io_data; // @[aes.scala 20:19:@2107.4]
  wire  encm_io_en; // @[aes.scala 20:19:@2107.4]
  wire  ke_clock; // @[aes.scala 22:18:@2113.4]
  wire  ke_reset; // @[aes.scala 22:18:@2113.4]
  wire [31:0] ke_io_sboxio_addr; // @[aes.scala 22:18:@2113.4]
  wire [31:0] ke_io_sboxio_data; // @[aes.scala 22:18:@2113.4]
  wire [3:0] ke_io_round; // @[aes.scala 22:18:@2113.4]
  wire [127:0] ke_io_data; // @[aes.scala 22:18:@2113.4]
  wire [127:0] ke_io_key; // @[aes.scala 22:18:@2113.4]
  wire [31:0] sb_io_addr; // @[aes.scala 23:18:@2116.4]
  wire [31:0] sb_io_data; // @[aes.scala 23:18:@2116.4]
  wire [127:0] sb_io_addr2; // @[aes.scala 23:18:@2116.4]
  wire [127:0] sb_io_data2; // @[aes.scala 23:18:@2116.4]
  wire  _T_18; // @[aes.scala 44:17:@2136.4]
  wire [127:0] _T_19; // @[aes.scala 51:19:@2138.4]
  wire [3:0] _T_20; // @[aes.scala 55:20:@2143.4]
  enc encm ( // @[aes.scala 20:19:@2107.4]
    .clock(encm_clock),
    .reset(encm_reset),
    .io_rkey(encm_io_rkey),
    .io_done(encm_io_done),
    .io_sio_addr2(encm_io_sio_addr2),
    .io_sio_data2(encm_io_sio_data2),
    .io_out(encm_io_out),
    .io_roundOut(encm_io_roundOut),
    .io_data(encm_io_data),
    .io_en(encm_io_en)
  );
  expander ke ( // @[aes.scala 22:18:@2113.4]
    .clock(ke_clock),
    .reset(ke_reset),
    .io_sboxio_addr(ke_io_sboxio_addr),
    .io_sboxio_data(ke_io_sboxio_data),
    .io_round(ke_io_round),
    .io_data(ke_io_data),
    .io_key(ke_io_key)
  );
  sbox sb ( // @[aes.scala 23:18:@2116.4]
    .io_addr(sb_io_addr),
    .io_data(sb_io_data),
    .io_addr2(sb_io_addr2),
    .io_data2(sb_io_data2)
  );
  assign _T_18 = io_en ? encm_io_done : 1'h0; // @[aes.scala 44:17:@2136.4]
  assign _T_19 = encm_io_out; // @[aes.scala 51:19:@2138.4]
  assign _T_20 = encm_io_roundOut; // @[aes.scala 55:20:@2143.4]
  assign io_result = _T_19;
  assign io_done = _T_18;
  assign encm_clock = clock;
  assign encm_reset = reset;
  assign encm_io_rkey = ke_io_data;
  assign encm_io_sio_data2 = sb_io_data2;
  assign encm_io_data = io_iData;
  assign encm_io_en = io_en;
  assign ke_clock = clock;
  assign ke_reset = reset;
  assign ke_io_sboxio_data = sb_io_data;
  assign ke_io_round = _T_20;
  assign ke_io_key = io_key;
  assign sb_io_addr = ke_io_sboxio_addr;
  assign sb_io_addr2 = encm_io_sio_addr2;
endmodule
module aesctr( // @[:@2149.2]
  input          clock, // @[:@2150.4]
  input          reset, // @[:@2151.4]
  input  [127:0] io_intVect, // @[:@2152.4]
  output         io_newR, // @[:@2152.4]
  output [127:0] io_out, // @[:@2152.4]
  input  [127:0] io_data, // @[:@2152.4]
  input          io_en, // @[:@2152.4]
  input  [127:0] io_key // @[:@2152.4]
);
  wire  aes_clock; // @[aesctr.scala 24:19:@2154.4]
  wire  aes_reset; // @[aesctr.scala 24:19:@2154.4]
  wire [127:0] aes_io_result; // @[aesctr.scala 24:19:@2154.4]
  wire [127:0] aes_io_iData; // @[aesctr.scala 24:19:@2154.4]
  wire [127:0] aes_io_key; // @[aesctr.scala 24:19:@2154.4]
  wire  aes_io_done; // @[aesctr.scala 24:19:@2154.4]
  wire  aes_io_en; // @[aesctr.scala 24:19:@2154.4]
  wire [127:0] _T_10; // @[aesctr.scala 35:44:@2162.4]
  wire [127:0] _T_12; // @[aesctr.scala 35:16:@2163.4]
  aes aes ( // @[aesctr.scala 24:19:@2154.4]
    .clock(aes_clock),
    .reset(aes_reset),
    .io_result(aes_io_result),
    .io_iData(aes_io_iData),
    .io_key(aes_io_key),
    .io_done(aes_io_done),
    .io_en(aes_io_en)
  );
  assign _T_10 = aes_io_result ^ io_data; // @[aesctr.scala 35:44:@2162.4]
  assign _T_12 = aes_io_done ? _T_10 : 128'h0; // @[aesctr.scala 35:16:@2163.4]
  assign io_newR = aes_io_done;
  assign io_out = _T_12;
  assign aes_clock = clock;
  assign aes_reset = reset;
  assign aes_io_iData = io_intVect;
  assign aes_io_key = io_key;
  assign aes_io_en = io_en;
endmodule
module g128Multiplay( // @[:@2166.2]
  input  [127:0] io_x, // @[:@2169.4]
  input  [127:0] io_y, // @[:@2169.4]
  output [127:0] io_out // @[:@2169.4]
);
  wire  _T_530; // @[G128Multiplay.scala 37:16:@2433.4]
  wire [127:0] Z_1; // @[G128Multiplay.scala 38:7:@2435.4]
  wire  _T_534; // @[G128Multiplay.scala 45:18:@2442.4]
  wire  _T_536; // @[G128Multiplay.scala 45:22:@2443.4]
  wire [127:0] _T_538; // @[G128Multiplay.scala 48:24:@2445.6]
  wire [127:0] _T_542; // @[G128Multiplay.scala 51:31:@2451.6]
  wire [127:0] V_1; // @[G128Multiplay.scala 46:7:@2444.4]
  wire  _T_544; // @[G128Multiplay.scala 37:16:@2455.4]
  wire [127:0] _T_547; // @[G128Multiplay.scala 40:24:@2458.6]
  wire [127:0] Z_2; // @[G128Multiplay.scala 38:7:@2457.4]
  wire  _T_548; // @[G128Multiplay.scala 45:18:@2464.4]
  wire  _T_550; // @[G128Multiplay.scala 45:22:@2465.4]
  wire [127:0] _T_552; // @[G128Multiplay.scala 48:24:@2467.6]
  wire [127:0] _T_556; // @[G128Multiplay.scala 51:31:@2473.6]
  wire [127:0] V_2; // @[G128Multiplay.scala 46:7:@2466.4]
  wire  _T_558; // @[G128Multiplay.scala 37:16:@2477.4]
  wire [127:0] _T_561; // @[G128Multiplay.scala 40:24:@2480.6]
  wire [127:0] Z_3; // @[G128Multiplay.scala 38:7:@2479.4]
  wire  _T_562; // @[G128Multiplay.scala 45:18:@2486.4]
  wire  _T_564; // @[G128Multiplay.scala 45:22:@2487.4]
  wire [127:0] _T_566; // @[G128Multiplay.scala 48:24:@2489.6]
  wire [127:0] _T_570; // @[G128Multiplay.scala 51:31:@2495.6]
  wire [127:0] V_3; // @[G128Multiplay.scala 46:7:@2488.4]
  wire  _T_572; // @[G128Multiplay.scala 37:16:@2499.4]
  wire [127:0] _T_575; // @[G128Multiplay.scala 40:24:@2502.6]
  wire [127:0] Z_4; // @[G128Multiplay.scala 38:7:@2501.4]
  wire  _T_576; // @[G128Multiplay.scala 45:18:@2508.4]
  wire  _T_578; // @[G128Multiplay.scala 45:22:@2509.4]
  wire [127:0] _T_580; // @[G128Multiplay.scala 48:24:@2511.6]
  wire [127:0] _T_584; // @[G128Multiplay.scala 51:31:@2517.6]
  wire [127:0] V_4; // @[G128Multiplay.scala 46:7:@2510.4]
  wire  _T_586; // @[G128Multiplay.scala 37:16:@2521.4]
  wire [127:0] _T_589; // @[G128Multiplay.scala 40:24:@2524.6]
  wire [127:0] Z_5; // @[G128Multiplay.scala 38:7:@2523.4]
  wire  _T_590; // @[G128Multiplay.scala 45:18:@2530.4]
  wire  _T_592; // @[G128Multiplay.scala 45:22:@2531.4]
  wire [127:0] _T_594; // @[G128Multiplay.scala 48:24:@2533.6]
  wire [127:0] _T_598; // @[G128Multiplay.scala 51:31:@2539.6]
  wire [127:0] V_5; // @[G128Multiplay.scala 46:7:@2532.4]
  wire  _T_600; // @[G128Multiplay.scala 37:16:@2543.4]
  wire [127:0] _T_603; // @[G128Multiplay.scala 40:24:@2546.6]
  wire [127:0] Z_6; // @[G128Multiplay.scala 38:7:@2545.4]
  wire  _T_604; // @[G128Multiplay.scala 45:18:@2552.4]
  wire  _T_606; // @[G128Multiplay.scala 45:22:@2553.4]
  wire [127:0] _T_608; // @[G128Multiplay.scala 48:24:@2555.6]
  wire [127:0] _T_612; // @[G128Multiplay.scala 51:31:@2561.6]
  wire [127:0] V_6; // @[G128Multiplay.scala 46:7:@2554.4]
  wire  _T_614; // @[G128Multiplay.scala 37:16:@2565.4]
  wire [127:0] _T_617; // @[G128Multiplay.scala 40:24:@2568.6]
  wire [127:0] Z_7; // @[G128Multiplay.scala 38:7:@2567.4]
  wire  _T_618; // @[G128Multiplay.scala 45:18:@2574.4]
  wire  _T_620; // @[G128Multiplay.scala 45:22:@2575.4]
  wire [127:0] _T_622; // @[G128Multiplay.scala 48:24:@2577.6]
  wire [127:0] _T_626; // @[G128Multiplay.scala 51:31:@2583.6]
  wire [127:0] V_7; // @[G128Multiplay.scala 46:7:@2576.4]
  wire  _T_628; // @[G128Multiplay.scala 37:16:@2587.4]
  wire [127:0] _T_631; // @[G128Multiplay.scala 40:24:@2590.6]
  wire [127:0] Z_8; // @[G128Multiplay.scala 38:7:@2589.4]
  wire  _T_632; // @[G128Multiplay.scala 45:18:@2596.4]
  wire  _T_634; // @[G128Multiplay.scala 45:22:@2597.4]
  wire [127:0] _T_636; // @[G128Multiplay.scala 48:24:@2599.6]
  wire [127:0] _T_640; // @[G128Multiplay.scala 51:31:@2605.6]
  wire [127:0] V_8; // @[G128Multiplay.scala 46:7:@2598.4]
  wire  _T_642; // @[G128Multiplay.scala 37:16:@2609.4]
  wire [127:0] _T_645; // @[G128Multiplay.scala 40:24:@2612.6]
  wire [127:0] Z_9; // @[G128Multiplay.scala 38:7:@2611.4]
  wire  _T_646; // @[G128Multiplay.scala 45:18:@2618.4]
  wire  _T_648; // @[G128Multiplay.scala 45:22:@2619.4]
  wire [127:0] _T_650; // @[G128Multiplay.scala 48:24:@2621.6]
  wire [127:0] _T_654; // @[G128Multiplay.scala 51:31:@2627.6]
  wire [127:0] V_9; // @[G128Multiplay.scala 46:7:@2620.4]
  wire  _T_656; // @[G128Multiplay.scala 37:16:@2631.4]
  wire [127:0] _T_659; // @[G128Multiplay.scala 40:24:@2634.6]
  wire [127:0] Z_10; // @[G128Multiplay.scala 38:7:@2633.4]
  wire  _T_660; // @[G128Multiplay.scala 45:18:@2640.4]
  wire  _T_662; // @[G128Multiplay.scala 45:22:@2641.4]
  wire [127:0] _T_664; // @[G128Multiplay.scala 48:24:@2643.6]
  wire [127:0] _T_668; // @[G128Multiplay.scala 51:31:@2649.6]
  wire [127:0] V_10; // @[G128Multiplay.scala 46:7:@2642.4]
  wire  _T_670; // @[G128Multiplay.scala 37:16:@2653.4]
  wire [127:0] _T_673; // @[G128Multiplay.scala 40:24:@2656.6]
  wire [127:0] Z_11; // @[G128Multiplay.scala 38:7:@2655.4]
  wire  _T_674; // @[G128Multiplay.scala 45:18:@2662.4]
  wire  _T_676; // @[G128Multiplay.scala 45:22:@2663.4]
  wire [127:0] _T_678; // @[G128Multiplay.scala 48:24:@2665.6]
  wire [127:0] _T_682; // @[G128Multiplay.scala 51:31:@2671.6]
  wire [127:0] V_11; // @[G128Multiplay.scala 46:7:@2664.4]
  wire  _T_684; // @[G128Multiplay.scala 37:16:@2675.4]
  wire [127:0] _T_687; // @[G128Multiplay.scala 40:24:@2678.6]
  wire [127:0] Z_12; // @[G128Multiplay.scala 38:7:@2677.4]
  wire  _T_688; // @[G128Multiplay.scala 45:18:@2684.4]
  wire  _T_690; // @[G128Multiplay.scala 45:22:@2685.4]
  wire [127:0] _T_692; // @[G128Multiplay.scala 48:24:@2687.6]
  wire [127:0] _T_696; // @[G128Multiplay.scala 51:31:@2693.6]
  wire [127:0] V_12; // @[G128Multiplay.scala 46:7:@2686.4]
  wire  _T_698; // @[G128Multiplay.scala 37:16:@2697.4]
  wire [127:0] _T_701; // @[G128Multiplay.scala 40:24:@2700.6]
  wire [127:0] Z_13; // @[G128Multiplay.scala 38:7:@2699.4]
  wire  _T_702; // @[G128Multiplay.scala 45:18:@2706.4]
  wire  _T_704; // @[G128Multiplay.scala 45:22:@2707.4]
  wire [127:0] _T_706; // @[G128Multiplay.scala 48:24:@2709.6]
  wire [127:0] _T_710; // @[G128Multiplay.scala 51:31:@2715.6]
  wire [127:0] V_13; // @[G128Multiplay.scala 46:7:@2708.4]
  wire  _T_712; // @[G128Multiplay.scala 37:16:@2719.4]
  wire [127:0] _T_715; // @[G128Multiplay.scala 40:24:@2722.6]
  wire [127:0] Z_14; // @[G128Multiplay.scala 38:7:@2721.4]
  wire  _T_716; // @[G128Multiplay.scala 45:18:@2728.4]
  wire  _T_718; // @[G128Multiplay.scala 45:22:@2729.4]
  wire [127:0] _T_720; // @[G128Multiplay.scala 48:24:@2731.6]
  wire [127:0] _T_724; // @[G128Multiplay.scala 51:31:@2737.6]
  wire [127:0] V_14; // @[G128Multiplay.scala 46:7:@2730.4]
  wire  _T_726; // @[G128Multiplay.scala 37:16:@2741.4]
  wire [127:0] _T_729; // @[G128Multiplay.scala 40:24:@2744.6]
  wire [127:0] Z_15; // @[G128Multiplay.scala 38:7:@2743.4]
  wire  _T_730; // @[G128Multiplay.scala 45:18:@2750.4]
  wire  _T_732; // @[G128Multiplay.scala 45:22:@2751.4]
  wire [127:0] _T_734; // @[G128Multiplay.scala 48:24:@2753.6]
  wire [127:0] _T_738; // @[G128Multiplay.scala 51:31:@2759.6]
  wire [127:0] V_15; // @[G128Multiplay.scala 46:7:@2752.4]
  wire  _T_740; // @[G128Multiplay.scala 37:16:@2763.4]
  wire [127:0] _T_743; // @[G128Multiplay.scala 40:24:@2766.6]
  wire [127:0] Z_16; // @[G128Multiplay.scala 38:7:@2765.4]
  wire  _T_744; // @[G128Multiplay.scala 45:18:@2772.4]
  wire  _T_746; // @[G128Multiplay.scala 45:22:@2773.4]
  wire [127:0] _T_748; // @[G128Multiplay.scala 48:24:@2775.6]
  wire [127:0] _T_752; // @[G128Multiplay.scala 51:31:@2781.6]
  wire [127:0] V_16; // @[G128Multiplay.scala 46:7:@2774.4]
  wire  _T_754; // @[G128Multiplay.scala 37:16:@2785.4]
  wire [127:0] _T_757; // @[G128Multiplay.scala 40:24:@2788.6]
  wire [127:0] Z_17; // @[G128Multiplay.scala 38:7:@2787.4]
  wire  _T_758; // @[G128Multiplay.scala 45:18:@2794.4]
  wire  _T_760; // @[G128Multiplay.scala 45:22:@2795.4]
  wire [127:0] _T_762; // @[G128Multiplay.scala 48:24:@2797.6]
  wire [127:0] _T_766; // @[G128Multiplay.scala 51:31:@2803.6]
  wire [127:0] V_17; // @[G128Multiplay.scala 46:7:@2796.4]
  wire  _T_768; // @[G128Multiplay.scala 37:16:@2807.4]
  wire [127:0] _T_771; // @[G128Multiplay.scala 40:24:@2810.6]
  wire [127:0] Z_18; // @[G128Multiplay.scala 38:7:@2809.4]
  wire  _T_772; // @[G128Multiplay.scala 45:18:@2816.4]
  wire  _T_774; // @[G128Multiplay.scala 45:22:@2817.4]
  wire [127:0] _T_776; // @[G128Multiplay.scala 48:24:@2819.6]
  wire [127:0] _T_780; // @[G128Multiplay.scala 51:31:@2825.6]
  wire [127:0] V_18; // @[G128Multiplay.scala 46:7:@2818.4]
  wire  _T_782; // @[G128Multiplay.scala 37:16:@2829.4]
  wire [127:0] _T_785; // @[G128Multiplay.scala 40:24:@2832.6]
  wire [127:0] Z_19; // @[G128Multiplay.scala 38:7:@2831.4]
  wire  _T_786; // @[G128Multiplay.scala 45:18:@2838.4]
  wire  _T_788; // @[G128Multiplay.scala 45:22:@2839.4]
  wire [127:0] _T_790; // @[G128Multiplay.scala 48:24:@2841.6]
  wire [127:0] _T_794; // @[G128Multiplay.scala 51:31:@2847.6]
  wire [127:0] V_19; // @[G128Multiplay.scala 46:7:@2840.4]
  wire  _T_796; // @[G128Multiplay.scala 37:16:@2851.4]
  wire [127:0] _T_799; // @[G128Multiplay.scala 40:24:@2854.6]
  wire [127:0] Z_20; // @[G128Multiplay.scala 38:7:@2853.4]
  wire  _T_800; // @[G128Multiplay.scala 45:18:@2860.4]
  wire  _T_802; // @[G128Multiplay.scala 45:22:@2861.4]
  wire [127:0] _T_804; // @[G128Multiplay.scala 48:24:@2863.6]
  wire [127:0] _T_808; // @[G128Multiplay.scala 51:31:@2869.6]
  wire [127:0] V_20; // @[G128Multiplay.scala 46:7:@2862.4]
  wire  _T_810; // @[G128Multiplay.scala 37:16:@2873.4]
  wire [127:0] _T_813; // @[G128Multiplay.scala 40:24:@2876.6]
  wire [127:0] Z_21; // @[G128Multiplay.scala 38:7:@2875.4]
  wire  _T_814; // @[G128Multiplay.scala 45:18:@2882.4]
  wire  _T_816; // @[G128Multiplay.scala 45:22:@2883.4]
  wire [127:0] _T_818; // @[G128Multiplay.scala 48:24:@2885.6]
  wire [127:0] _T_822; // @[G128Multiplay.scala 51:31:@2891.6]
  wire [127:0] V_21; // @[G128Multiplay.scala 46:7:@2884.4]
  wire  _T_824; // @[G128Multiplay.scala 37:16:@2895.4]
  wire [127:0] _T_827; // @[G128Multiplay.scala 40:24:@2898.6]
  wire [127:0] Z_22; // @[G128Multiplay.scala 38:7:@2897.4]
  wire  _T_828; // @[G128Multiplay.scala 45:18:@2904.4]
  wire  _T_830; // @[G128Multiplay.scala 45:22:@2905.4]
  wire [127:0] _T_832; // @[G128Multiplay.scala 48:24:@2907.6]
  wire [127:0] _T_836; // @[G128Multiplay.scala 51:31:@2913.6]
  wire [127:0] V_22; // @[G128Multiplay.scala 46:7:@2906.4]
  wire  _T_838; // @[G128Multiplay.scala 37:16:@2917.4]
  wire [127:0] _T_841; // @[G128Multiplay.scala 40:24:@2920.6]
  wire [127:0] Z_23; // @[G128Multiplay.scala 38:7:@2919.4]
  wire  _T_842; // @[G128Multiplay.scala 45:18:@2926.4]
  wire  _T_844; // @[G128Multiplay.scala 45:22:@2927.4]
  wire [127:0] _T_846; // @[G128Multiplay.scala 48:24:@2929.6]
  wire [127:0] _T_850; // @[G128Multiplay.scala 51:31:@2935.6]
  wire [127:0] V_23; // @[G128Multiplay.scala 46:7:@2928.4]
  wire  _T_852; // @[G128Multiplay.scala 37:16:@2939.4]
  wire [127:0] _T_855; // @[G128Multiplay.scala 40:24:@2942.6]
  wire [127:0] Z_24; // @[G128Multiplay.scala 38:7:@2941.4]
  wire  _T_856; // @[G128Multiplay.scala 45:18:@2948.4]
  wire  _T_858; // @[G128Multiplay.scala 45:22:@2949.4]
  wire [127:0] _T_860; // @[G128Multiplay.scala 48:24:@2951.6]
  wire [127:0] _T_864; // @[G128Multiplay.scala 51:31:@2957.6]
  wire [127:0] V_24; // @[G128Multiplay.scala 46:7:@2950.4]
  wire  _T_866; // @[G128Multiplay.scala 37:16:@2961.4]
  wire [127:0] _T_869; // @[G128Multiplay.scala 40:24:@2964.6]
  wire [127:0] Z_25; // @[G128Multiplay.scala 38:7:@2963.4]
  wire  _T_870; // @[G128Multiplay.scala 45:18:@2970.4]
  wire  _T_872; // @[G128Multiplay.scala 45:22:@2971.4]
  wire [127:0] _T_874; // @[G128Multiplay.scala 48:24:@2973.6]
  wire [127:0] _T_878; // @[G128Multiplay.scala 51:31:@2979.6]
  wire [127:0] V_25; // @[G128Multiplay.scala 46:7:@2972.4]
  wire  _T_880; // @[G128Multiplay.scala 37:16:@2983.4]
  wire [127:0] _T_883; // @[G128Multiplay.scala 40:24:@2986.6]
  wire [127:0] Z_26; // @[G128Multiplay.scala 38:7:@2985.4]
  wire  _T_884; // @[G128Multiplay.scala 45:18:@2992.4]
  wire  _T_886; // @[G128Multiplay.scala 45:22:@2993.4]
  wire [127:0] _T_888; // @[G128Multiplay.scala 48:24:@2995.6]
  wire [127:0] _T_892; // @[G128Multiplay.scala 51:31:@3001.6]
  wire [127:0] V_26; // @[G128Multiplay.scala 46:7:@2994.4]
  wire  _T_894; // @[G128Multiplay.scala 37:16:@3005.4]
  wire [127:0] _T_897; // @[G128Multiplay.scala 40:24:@3008.6]
  wire [127:0] Z_27; // @[G128Multiplay.scala 38:7:@3007.4]
  wire  _T_898; // @[G128Multiplay.scala 45:18:@3014.4]
  wire  _T_900; // @[G128Multiplay.scala 45:22:@3015.4]
  wire [127:0] _T_902; // @[G128Multiplay.scala 48:24:@3017.6]
  wire [127:0] _T_906; // @[G128Multiplay.scala 51:31:@3023.6]
  wire [127:0] V_27; // @[G128Multiplay.scala 46:7:@3016.4]
  wire  _T_908; // @[G128Multiplay.scala 37:16:@3027.4]
  wire [127:0] _T_911; // @[G128Multiplay.scala 40:24:@3030.6]
  wire [127:0] Z_28; // @[G128Multiplay.scala 38:7:@3029.4]
  wire  _T_912; // @[G128Multiplay.scala 45:18:@3036.4]
  wire  _T_914; // @[G128Multiplay.scala 45:22:@3037.4]
  wire [127:0] _T_916; // @[G128Multiplay.scala 48:24:@3039.6]
  wire [127:0] _T_920; // @[G128Multiplay.scala 51:31:@3045.6]
  wire [127:0] V_28; // @[G128Multiplay.scala 46:7:@3038.4]
  wire  _T_922; // @[G128Multiplay.scala 37:16:@3049.4]
  wire [127:0] _T_925; // @[G128Multiplay.scala 40:24:@3052.6]
  wire [127:0] Z_29; // @[G128Multiplay.scala 38:7:@3051.4]
  wire  _T_926; // @[G128Multiplay.scala 45:18:@3058.4]
  wire  _T_928; // @[G128Multiplay.scala 45:22:@3059.4]
  wire [127:0] _T_930; // @[G128Multiplay.scala 48:24:@3061.6]
  wire [127:0] _T_934; // @[G128Multiplay.scala 51:31:@3067.6]
  wire [127:0] V_29; // @[G128Multiplay.scala 46:7:@3060.4]
  wire  _T_936; // @[G128Multiplay.scala 37:16:@3071.4]
  wire [127:0] _T_939; // @[G128Multiplay.scala 40:24:@3074.6]
  wire [127:0] Z_30; // @[G128Multiplay.scala 38:7:@3073.4]
  wire  _T_940; // @[G128Multiplay.scala 45:18:@3080.4]
  wire  _T_942; // @[G128Multiplay.scala 45:22:@3081.4]
  wire [127:0] _T_944; // @[G128Multiplay.scala 48:24:@3083.6]
  wire [127:0] _T_948; // @[G128Multiplay.scala 51:31:@3089.6]
  wire [127:0] V_30; // @[G128Multiplay.scala 46:7:@3082.4]
  wire  _T_950; // @[G128Multiplay.scala 37:16:@3093.4]
  wire [127:0] _T_953; // @[G128Multiplay.scala 40:24:@3096.6]
  wire [127:0] Z_31; // @[G128Multiplay.scala 38:7:@3095.4]
  wire  _T_954; // @[G128Multiplay.scala 45:18:@3102.4]
  wire  _T_956; // @[G128Multiplay.scala 45:22:@3103.4]
  wire [127:0] _T_958; // @[G128Multiplay.scala 48:24:@3105.6]
  wire [127:0] _T_962; // @[G128Multiplay.scala 51:31:@3111.6]
  wire [127:0] V_31; // @[G128Multiplay.scala 46:7:@3104.4]
  wire  _T_964; // @[G128Multiplay.scala 37:16:@3115.4]
  wire [127:0] _T_967; // @[G128Multiplay.scala 40:24:@3118.6]
  wire [127:0] Z_32; // @[G128Multiplay.scala 38:7:@3117.4]
  wire  _T_968; // @[G128Multiplay.scala 45:18:@3124.4]
  wire  _T_970; // @[G128Multiplay.scala 45:22:@3125.4]
  wire [127:0] _T_972; // @[G128Multiplay.scala 48:24:@3127.6]
  wire [127:0] _T_976; // @[G128Multiplay.scala 51:31:@3133.6]
  wire [127:0] V_32; // @[G128Multiplay.scala 46:7:@3126.4]
  wire  _T_978; // @[G128Multiplay.scala 37:16:@3137.4]
  wire [127:0] _T_981; // @[G128Multiplay.scala 40:24:@3140.6]
  wire [127:0] Z_33; // @[G128Multiplay.scala 38:7:@3139.4]
  wire  _T_982; // @[G128Multiplay.scala 45:18:@3146.4]
  wire  _T_984; // @[G128Multiplay.scala 45:22:@3147.4]
  wire [127:0] _T_986; // @[G128Multiplay.scala 48:24:@3149.6]
  wire [127:0] _T_990; // @[G128Multiplay.scala 51:31:@3155.6]
  wire [127:0] V_33; // @[G128Multiplay.scala 46:7:@3148.4]
  wire  _T_992; // @[G128Multiplay.scala 37:16:@3159.4]
  wire [127:0] _T_995; // @[G128Multiplay.scala 40:24:@3162.6]
  wire [127:0] Z_34; // @[G128Multiplay.scala 38:7:@3161.4]
  wire  _T_996; // @[G128Multiplay.scala 45:18:@3168.4]
  wire  _T_998; // @[G128Multiplay.scala 45:22:@3169.4]
  wire [127:0] _T_1000; // @[G128Multiplay.scala 48:24:@3171.6]
  wire [127:0] _T_1004; // @[G128Multiplay.scala 51:31:@3177.6]
  wire [127:0] V_34; // @[G128Multiplay.scala 46:7:@3170.4]
  wire  _T_1006; // @[G128Multiplay.scala 37:16:@3181.4]
  wire [127:0] _T_1009; // @[G128Multiplay.scala 40:24:@3184.6]
  wire [127:0] Z_35; // @[G128Multiplay.scala 38:7:@3183.4]
  wire  _T_1010; // @[G128Multiplay.scala 45:18:@3190.4]
  wire  _T_1012; // @[G128Multiplay.scala 45:22:@3191.4]
  wire [127:0] _T_1014; // @[G128Multiplay.scala 48:24:@3193.6]
  wire [127:0] _T_1018; // @[G128Multiplay.scala 51:31:@3199.6]
  wire [127:0] V_35; // @[G128Multiplay.scala 46:7:@3192.4]
  wire  _T_1020; // @[G128Multiplay.scala 37:16:@3203.4]
  wire [127:0] _T_1023; // @[G128Multiplay.scala 40:24:@3206.6]
  wire [127:0] Z_36; // @[G128Multiplay.scala 38:7:@3205.4]
  wire  _T_1024; // @[G128Multiplay.scala 45:18:@3212.4]
  wire  _T_1026; // @[G128Multiplay.scala 45:22:@3213.4]
  wire [127:0] _T_1028; // @[G128Multiplay.scala 48:24:@3215.6]
  wire [127:0] _T_1032; // @[G128Multiplay.scala 51:31:@3221.6]
  wire [127:0] V_36; // @[G128Multiplay.scala 46:7:@3214.4]
  wire  _T_1034; // @[G128Multiplay.scala 37:16:@3225.4]
  wire [127:0] _T_1037; // @[G128Multiplay.scala 40:24:@3228.6]
  wire [127:0] Z_37; // @[G128Multiplay.scala 38:7:@3227.4]
  wire  _T_1038; // @[G128Multiplay.scala 45:18:@3234.4]
  wire  _T_1040; // @[G128Multiplay.scala 45:22:@3235.4]
  wire [127:0] _T_1042; // @[G128Multiplay.scala 48:24:@3237.6]
  wire [127:0] _T_1046; // @[G128Multiplay.scala 51:31:@3243.6]
  wire [127:0] V_37; // @[G128Multiplay.scala 46:7:@3236.4]
  wire  _T_1048; // @[G128Multiplay.scala 37:16:@3247.4]
  wire [127:0] _T_1051; // @[G128Multiplay.scala 40:24:@3250.6]
  wire [127:0] Z_38; // @[G128Multiplay.scala 38:7:@3249.4]
  wire  _T_1052; // @[G128Multiplay.scala 45:18:@3256.4]
  wire  _T_1054; // @[G128Multiplay.scala 45:22:@3257.4]
  wire [127:0] _T_1056; // @[G128Multiplay.scala 48:24:@3259.6]
  wire [127:0] _T_1060; // @[G128Multiplay.scala 51:31:@3265.6]
  wire [127:0] V_38; // @[G128Multiplay.scala 46:7:@3258.4]
  wire  _T_1062; // @[G128Multiplay.scala 37:16:@3269.4]
  wire [127:0] _T_1065; // @[G128Multiplay.scala 40:24:@3272.6]
  wire [127:0] Z_39; // @[G128Multiplay.scala 38:7:@3271.4]
  wire  _T_1066; // @[G128Multiplay.scala 45:18:@3278.4]
  wire  _T_1068; // @[G128Multiplay.scala 45:22:@3279.4]
  wire [127:0] _T_1070; // @[G128Multiplay.scala 48:24:@3281.6]
  wire [127:0] _T_1074; // @[G128Multiplay.scala 51:31:@3287.6]
  wire [127:0] V_39; // @[G128Multiplay.scala 46:7:@3280.4]
  wire  _T_1076; // @[G128Multiplay.scala 37:16:@3291.4]
  wire [127:0] _T_1079; // @[G128Multiplay.scala 40:24:@3294.6]
  wire [127:0] Z_40; // @[G128Multiplay.scala 38:7:@3293.4]
  wire  _T_1080; // @[G128Multiplay.scala 45:18:@3300.4]
  wire  _T_1082; // @[G128Multiplay.scala 45:22:@3301.4]
  wire [127:0] _T_1084; // @[G128Multiplay.scala 48:24:@3303.6]
  wire [127:0] _T_1088; // @[G128Multiplay.scala 51:31:@3309.6]
  wire [127:0] V_40; // @[G128Multiplay.scala 46:7:@3302.4]
  wire  _T_1090; // @[G128Multiplay.scala 37:16:@3313.4]
  wire [127:0] _T_1093; // @[G128Multiplay.scala 40:24:@3316.6]
  wire [127:0] Z_41; // @[G128Multiplay.scala 38:7:@3315.4]
  wire  _T_1094; // @[G128Multiplay.scala 45:18:@3322.4]
  wire  _T_1096; // @[G128Multiplay.scala 45:22:@3323.4]
  wire [127:0] _T_1098; // @[G128Multiplay.scala 48:24:@3325.6]
  wire [127:0] _T_1102; // @[G128Multiplay.scala 51:31:@3331.6]
  wire [127:0] V_41; // @[G128Multiplay.scala 46:7:@3324.4]
  wire  _T_1104; // @[G128Multiplay.scala 37:16:@3335.4]
  wire [127:0] _T_1107; // @[G128Multiplay.scala 40:24:@3338.6]
  wire [127:0] Z_42; // @[G128Multiplay.scala 38:7:@3337.4]
  wire  _T_1108; // @[G128Multiplay.scala 45:18:@3344.4]
  wire  _T_1110; // @[G128Multiplay.scala 45:22:@3345.4]
  wire [127:0] _T_1112; // @[G128Multiplay.scala 48:24:@3347.6]
  wire [127:0] _T_1116; // @[G128Multiplay.scala 51:31:@3353.6]
  wire [127:0] V_42; // @[G128Multiplay.scala 46:7:@3346.4]
  wire  _T_1118; // @[G128Multiplay.scala 37:16:@3357.4]
  wire [127:0] _T_1121; // @[G128Multiplay.scala 40:24:@3360.6]
  wire [127:0] Z_43; // @[G128Multiplay.scala 38:7:@3359.4]
  wire  _T_1122; // @[G128Multiplay.scala 45:18:@3366.4]
  wire  _T_1124; // @[G128Multiplay.scala 45:22:@3367.4]
  wire [127:0] _T_1126; // @[G128Multiplay.scala 48:24:@3369.6]
  wire [127:0] _T_1130; // @[G128Multiplay.scala 51:31:@3375.6]
  wire [127:0] V_43; // @[G128Multiplay.scala 46:7:@3368.4]
  wire  _T_1132; // @[G128Multiplay.scala 37:16:@3379.4]
  wire [127:0] _T_1135; // @[G128Multiplay.scala 40:24:@3382.6]
  wire [127:0] Z_44; // @[G128Multiplay.scala 38:7:@3381.4]
  wire  _T_1136; // @[G128Multiplay.scala 45:18:@3388.4]
  wire  _T_1138; // @[G128Multiplay.scala 45:22:@3389.4]
  wire [127:0] _T_1140; // @[G128Multiplay.scala 48:24:@3391.6]
  wire [127:0] _T_1144; // @[G128Multiplay.scala 51:31:@3397.6]
  wire [127:0] V_44; // @[G128Multiplay.scala 46:7:@3390.4]
  wire  _T_1146; // @[G128Multiplay.scala 37:16:@3401.4]
  wire [127:0] _T_1149; // @[G128Multiplay.scala 40:24:@3404.6]
  wire [127:0] Z_45; // @[G128Multiplay.scala 38:7:@3403.4]
  wire  _T_1150; // @[G128Multiplay.scala 45:18:@3410.4]
  wire  _T_1152; // @[G128Multiplay.scala 45:22:@3411.4]
  wire [127:0] _T_1154; // @[G128Multiplay.scala 48:24:@3413.6]
  wire [127:0] _T_1158; // @[G128Multiplay.scala 51:31:@3419.6]
  wire [127:0] V_45; // @[G128Multiplay.scala 46:7:@3412.4]
  wire  _T_1160; // @[G128Multiplay.scala 37:16:@3423.4]
  wire [127:0] _T_1163; // @[G128Multiplay.scala 40:24:@3426.6]
  wire [127:0] Z_46; // @[G128Multiplay.scala 38:7:@3425.4]
  wire  _T_1164; // @[G128Multiplay.scala 45:18:@3432.4]
  wire  _T_1166; // @[G128Multiplay.scala 45:22:@3433.4]
  wire [127:0] _T_1168; // @[G128Multiplay.scala 48:24:@3435.6]
  wire [127:0] _T_1172; // @[G128Multiplay.scala 51:31:@3441.6]
  wire [127:0] V_46; // @[G128Multiplay.scala 46:7:@3434.4]
  wire  _T_1174; // @[G128Multiplay.scala 37:16:@3445.4]
  wire [127:0] _T_1177; // @[G128Multiplay.scala 40:24:@3448.6]
  wire [127:0] Z_47; // @[G128Multiplay.scala 38:7:@3447.4]
  wire  _T_1178; // @[G128Multiplay.scala 45:18:@3454.4]
  wire  _T_1180; // @[G128Multiplay.scala 45:22:@3455.4]
  wire [127:0] _T_1182; // @[G128Multiplay.scala 48:24:@3457.6]
  wire [127:0] _T_1186; // @[G128Multiplay.scala 51:31:@3463.6]
  wire [127:0] V_47; // @[G128Multiplay.scala 46:7:@3456.4]
  wire  _T_1188; // @[G128Multiplay.scala 37:16:@3467.4]
  wire [127:0] _T_1191; // @[G128Multiplay.scala 40:24:@3470.6]
  wire [127:0] Z_48; // @[G128Multiplay.scala 38:7:@3469.4]
  wire  _T_1192; // @[G128Multiplay.scala 45:18:@3476.4]
  wire  _T_1194; // @[G128Multiplay.scala 45:22:@3477.4]
  wire [127:0] _T_1196; // @[G128Multiplay.scala 48:24:@3479.6]
  wire [127:0] _T_1200; // @[G128Multiplay.scala 51:31:@3485.6]
  wire [127:0] V_48; // @[G128Multiplay.scala 46:7:@3478.4]
  wire  _T_1202; // @[G128Multiplay.scala 37:16:@3489.4]
  wire [127:0] _T_1205; // @[G128Multiplay.scala 40:24:@3492.6]
  wire [127:0] Z_49; // @[G128Multiplay.scala 38:7:@3491.4]
  wire  _T_1206; // @[G128Multiplay.scala 45:18:@3498.4]
  wire  _T_1208; // @[G128Multiplay.scala 45:22:@3499.4]
  wire [127:0] _T_1210; // @[G128Multiplay.scala 48:24:@3501.6]
  wire [127:0] _T_1214; // @[G128Multiplay.scala 51:31:@3507.6]
  wire [127:0] V_49; // @[G128Multiplay.scala 46:7:@3500.4]
  wire  _T_1216; // @[G128Multiplay.scala 37:16:@3511.4]
  wire [127:0] _T_1219; // @[G128Multiplay.scala 40:24:@3514.6]
  wire [127:0] Z_50; // @[G128Multiplay.scala 38:7:@3513.4]
  wire  _T_1220; // @[G128Multiplay.scala 45:18:@3520.4]
  wire  _T_1222; // @[G128Multiplay.scala 45:22:@3521.4]
  wire [127:0] _T_1224; // @[G128Multiplay.scala 48:24:@3523.6]
  wire [127:0] _T_1228; // @[G128Multiplay.scala 51:31:@3529.6]
  wire [127:0] V_50; // @[G128Multiplay.scala 46:7:@3522.4]
  wire  _T_1230; // @[G128Multiplay.scala 37:16:@3533.4]
  wire [127:0] _T_1233; // @[G128Multiplay.scala 40:24:@3536.6]
  wire [127:0] Z_51; // @[G128Multiplay.scala 38:7:@3535.4]
  wire  _T_1234; // @[G128Multiplay.scala 45:18:@3542.4]
  wire  _T_1236; // @[G128Multiplay.scala 45:22:@3543.4]
  wire [127:0] _T_1238; // @[G128Multiplay.scala 48:24:@3545.6]
  wire [127:0] _T_1242; // @[G128Multiplay.scala 51:31:@3551.6]
  wire [127:0] V_51; // @[G128Multiplay.scala 46:7:@3544.4]
  wire  _T_1244; // @[G128Multiplay.scala 37:16:@3555.4]
  wire [127:0] _T_1247; // @[G128Multiplay.scala 40:24:@3558.6]
  wire [127:0] Z_52; // @[G128Multiplay.scala 38:7:@3557.4]
  wire  _T_1248; // @[G128Multiplay.scala 45:18:@3564.4]
  wire  _T_1250; // @[G128Multiplay.scala 45:22:@3565.4]
  wire [127:0] _T_1252; // @[G128Multiplay.scala 48:24:@3567.6]
  wire [127:0] _T_1256; // @[G128Multiplay.scala 51:31:@3573.6]
  wire [127:0] V_52; // @[G128Multiplay.scala 46:7:@3566.4]
  wire  _T_1258; // @[G128Multiplay.scala 37:16:@3577.4]
  wire [127:0] _T_1261; // @[G128Multiplay.scala 40:24:@3580.6]
  wire [127:0] Z_53; // @[G128Multiplay.scala 38:7:@3579.4]
  wire  _T_1262; // @[G128Multiplay.scala 45:18:@3586.4]
  wire  _T_1264; // @[G128Multiplay.scala 45:22:@3587.4]
  wire [127:0] _T_1266; // @[G128Multiplay.scala 48:24:@3589.6]
  wire [127:0] _T_1270; // @[G128Multiplay.scala 51:31:@3595.6]
  wire [127:0] V_53; // @[G128Multiplay.scala 46:7:@3588.4]
  wire  _T_1272; // @[G128Multiplay.scala 37:16:@3599.4]
  wire [127:0] _T_1275; // @[G128Multiplay.scala 40:24:@3602.6]
  wire [127:0] Z_54; // @[G128Multiplay.scala 38:7:@3601.4]
  wire  _T_1276; // @[G128Multiplay.scala 45:18:@3608.4]
  wire  _T_1278; // @[G128Multiplay.scala 45:22:@3609.4]
  wire [127:0] _T_1280; // @[G128Multiplay.scala 48:24:@3611.6]
  wire [127:0] _T_1284; // @[G128Multiplay.scala 51:31:@3617.6]
  wire [127:0] V_54; // @[G128Multiplay.scala 46:7:@3610.4]
  wire  _T_1286; // @[G128Multiplay.scala 37:16:@3621.4]
  wire [127:0] _T_1289; // @[G128Multiplay.scala 40:24:@3624.6]
  wire [127:0] Z_55; // @[G128Multiplay.scala 38:7:@3623.4]
  wire  _T_1290; // @[G128Multiplay.scala 45:18:@3630.4]
  wire  _T_1292; // @[G128Multiplay.scala 45:22:@3631.4]
  wire [127:0] _T_1294; // @[G128Multiplay.scala 48:24:@3633.6]
  wire [127:0] _T_1298; // @[G128Multiplay.scala 51:31:@3639.6]
  wire [127:0] V_55; // @[G128Multiplay.scala 46:7:@3632.4]
  wire  _T_1300; // @[G128Multiplay.scala 37:16:@3643.4]
  wire [127:0] _T_1303; // @[G128Multiplay.scala 40:24:@3646.6]
  wire [127:0] Z_56; // @[G128Multiplay.scala 38:7:@3645.4]
  wire  _T_1304; // @[G128Multiplay.scala 45:18:@3652.4]
  wire  _T_1306; // @[G128Multiplay.scala 45:22:@3653.4]
  wire [127:0] _T_1308; // @[G128Multiplay.scala 48:24:@3655.6]
  wire [127:0] _T_1312; // @[G128Multiplay.scala 51:31:@3661.6]
  wire [127:0] V_56; // @[G128Multiplay.scala 46:7:@3654.4]
  wire  _T_1314; // @[G128Multiplay.scala 37:16:@3665.4]
  wire [127:0] _T_1317; // @[G128Multiplay.scala 40:24:@3668.6]
  wire [127:0] Z_57; // @[G128Multiplay.scala 38:7:@3667.4]
  wire  _T_1318; // @[G128Multiplay.scala 45:18:@3674.4]
  wire  _T_1320; // @[G128Multiplay.scala 45:22:@3675.4]
  wire [127:0] _T_1322; // @[G128Multiplay.scala 48:24:@3677.6]
  wire [127:0] _T_1326; // @[G128Multiplay.scala 51:31:@3683.6]
  wire [127:0] V_57; // @[G128Multiplay.scala 46:7:@3676.4]
  wire  _T_1328; // @[G128Multiplay.scala 37:16:@3687.4]
  wire [127:0] _T_1331; // @[G128Multiplay.scala 40:24:@3690.6]
  wire [127:0] Z_58; // @[G128Multiplay.scala 38:7:@3689.4]
  wire  _T_1332; // @[G128Multiplay.scala 45:18:@3696.4]
  wire  _T_1334; // @[G128Multiplay.scala 45:22:@3697.4]
  wire [127:0] _T_1336; // @[G128Multiplay.scala 48:24:@3699.6]
  wire [127:0] _T_1340; // @[G128Multiplay.scala 51:31:@3705.6]
  wire [127:0] V_58; // @[G128Multiplay.scala 46:7:@3698.4]
  wire  _T_1342; // @[G128Multiplay.scala 37:16:@3709.4]
  wire [127:0] _T_1345; // @[G128Multiplay.scala 40:24:@3712.6]
  wire [127:0] Z_59; // @[G128Multiplay.scala 38:7:@3711.4]
  wire  _T_1346; // @[G128Multiplay.scala 45:18:@3718.4]
  wire  _T_1348; // @[G128Multiplay.scala 45:22:@3719.4]
  wire [127:0] _T_1350; // @[G128Multiplay.scala 48:24:@3721.6]
  wire [127:0] _T_1354; // @[G128Multiplay.scala 51:31:@3727.6]
  wire [127:0] V_59; // @[G128Multiplay.scala 46:7:@3720.4]
  wire  _T_1356; // @[G128Multiplay.scala 37:16:@3731.4]
  wire [127:0] _T_1359; // @[G128Multiplay.scala 40:24:@3734.6]
  wire [127:0] Z_60; // @[G128Multiplay.scala 38:7:@3733.4]
  wire  _T_1360; // @[G128Multiplay.scala 45:18:@3740.4]
  wire  _T_1362; // @[G128Multiplay.scala 45:22:@3741.4]
  wire [127:0] _T_1364; // @[G128Multiplay.scala 48:24:@3743.6]
  wire [127:0] _T_1368; // @[G128Multiplay.scala 51:31:@3749.6]
  wire [127:0] V_60; // @[G128Multiplay.scala 46:7:@3742.4]
  wire  _T_1370; // @[G128Multiplay.scala 37:16:@3753.4]
  wire [127:0] _T_1373; // @[G128Multiplay.scala 40:24:@3756.6]
  wire [127:0] Z_61; // @[G128Multiplay.scala 38:7:@3755.4]
  wire  _T_1374; // @[G128Multiplay.scala 45:18:@3762.4]
  wire  _T_1376; // @[G128Multiplay.scala 45:22:@3763.4]
  wire [127:0] _T_1378; // @[G128Multiplay.scala 48:24:@3765.6]
  wire [127:0] _T_1382; // @[G128Multiplay.scala 51:31:@3771.6]
  wire [127:0] V_61; // @[G128Multiplay.scala 46:7:@3764.4]
  wire  _T_1384; // @[G128Multiplay.scala 37:16:@3775.4]
  wire [127:0] _T_1387; // @[G128Multiplay.scala 40:24:@3778.6]
  wire [127:0] Z_62; // @[G128Multiplay.scala 38:7:@3777.4]
  wire  _T_1388; // @[G128Multiplay.scala 45:18:@3784.4]
  wire  _T_1390; // @[G128Multiplay.scala 45:22:@3785.4]
  wire [127:0] _T_1392; // @[G128Multiplay.scala 48:24:@3787.6]
  wire [127:0] _T_1396; // @[G128Multiplay.scala 51:31:@3793.6]
  wire [127:0] V_62; // @[G128Multiplay.scala 46:7:@3786.4]
  wire  _T_1398; // @[G128Multiplay.scala 37:16:@3797.4]
  wire [127:0] _T_1401; // @[G128Multiplay.scala 40:24:@3800.6]
  wire [127:0] Z_63; // @[G128Multiplay.scala 38:7:@3799.4]
  wire  _T_1402; // @[G128Multiplay.scala 45:18:@3806.4]
  wire  _T_1404; // @[G128Multiplay.scala 45:22:@3807.4]
  wire [127:0] _T_1406; // @[G128Multiplay.scala 48:24:@3809.6]
  wire [127:0] _T_1410; // @[G128Multiplay.scala 51:31:@3815.6]
  wire [127:0] V_63; // @[G128Multiplay.scala 46:7:@3808.4]
  wire  _T_1412; // @[G128Multiplay.scala 37:16:@3819.4]
  wire [127:0] _T_1415; // @[G128Multiplay.scala 40:24:@3822.6]
  wire [127:0] Z_64; // @[G128Multiplay.scala 38:7:@3821.4]
  wire  _T_1416; // @[G128Multiplay.scala 45:18:@3828.4]
  wire  _T_1418; // @[G128Multiplay.scala 45:22:@3829.4]
  wire [127:0] _T_1420; // @[G128Multiplay.scala 48:24:@3831.6]
  wire [127:0] _T_1424; // @[G128Multiplay.scala 51:31:@3837.6]
  wire [127:0] V_64; // @[G128Multiplay.scala 46:7:@3830.4]
  wire  _T_1426; // @[G128Multiplay.scala 37:16:@3841.4]
  wire [127:0] _T_1429; // @[G128Multiplay.scala 40:24:@3844.6]
  wire [127:0] Z_65; // @[G128Multiplay.scala 38:7:@3843.4]
  wire  _T_1430; // @[G128Multiplay.scala 45:18:@3850.4]
  wire  _T_1432; // @[G128Multiplay.scala 45:22:@3851.4]
  wire [127:0] _T_1434; // @[G128Multiplay.scala 48:24:@3853.6]
  wire [127:0] _T_1438; // @[G128Multiplay.scala 51:31:@3859.6]
  wire [127:0] V_65; // @[G128Multiplay.scala 46:7:@3852.4]
  wire  _T_1440; // @[G128Multiplay.scala 37:16:@3863.4]
  wire [127:0] _T_1443; // @[G128Multiplay.scala 40:24:@3866.6]
  wire [127:0] Z_66; // @[G128Multiplay.scala 38:7:@3865.4]
  wire  _T_1444; // @[G128Multiplay.scala 45:18:@3872.4]
  wire  _T_1446; // @[G128Multiplay.scala 45:22:@3873.4]
  wire [127:0] _T_1448; // @[G128Multiplay.scala 48:24:@3875.6]
  wire [127:0] _T_1452; // @[G128Multiplay.scala 51:31:@3881.6]
  wire [127:0] V_66; // @[G128Multiplay.scala 46:7:@3874.4]
  wire  _T_1454; // @[G128Multiplay.scala 37:16:@3885.4]
  wire [127:0] _T_1457; // @[G128Multiplay.scala 40:24:@3888.6]
  wire [127:0] Z_67; // @[G128Multiplay.scala 38:7:@3887.4]
  wire  _T_1458; // @[G128Multiplay.scala 45:18:@3894.4]
  wire  _T_1460; // @[G128Multiplay.scala 45:22:@3895.4]
  wire [127:0] _T_1462; // @[G128Multiplay.scala 48:24:@3897.6]
  wire [127:0] _T_1466; // @[G128Multiplay.scala 51:31:@3903.6]
  wire [127:0] V_67; // @[G128Multiplay.scala 46:7:@3896.4]
  wire  _T_1468; // @[G128Multiplay.scala 37:16:@3907.4]
  wire [127:0] _T_1471; // @[G128Multiplay.scala 40:24:@3910.6]
  wire [127:0] Z_68; // @[G128Multiplay.scala 38:7:@3909.4]
  wire  _T_1472; // @[G128Multiplay.scala 45:18:@3916.4]
  wire  _T_1474; // @[G128Multiplay.scala 45:22:@3917.4]
  wire [127:0] _T_1476; // @[G128Multiplay.scala 48:24:@3919.6]
  wire [127:0] _T_1480; // @[G128Multiplay.scala 51:31:@3925.6]
  wire [127:0] V_68; // @[G128Multiplay.scala 46:7:@3918.4]
  wire  _T_1482; // @[G128Multiplay.scala 37:16:@3929.4]
  wire [127:0] _T_1485; // @[G128Multiplay.scala 40:24:@3932.6]
  wire [127:0] Z_69; // @[G128Multiplay.scala 38:7:@3931.4]
  wire  _T_1486; // @[G128Multiplay.scala 45:18:@3938.4]
  wire  _T_1488; // @[G128Multiplay.scala 45:22:@3939.4]
  wire [127:0] _T_1490; // @[G128Multiplay.scala 48:24:@3941.6]
  wire [127:0] _T_1494; // @[G128Multiplay.scala 51:31:@3947.6]
  wire [127:0] V_69; // @[G128Multiplay.scala 46:7:@3940.4]
  wire  _T_1496; // @[G128Multiplay.scala 37:16:@3951.4]
  wire [127:0] _T_1499; // @[G128Multiplay.scala 40:24:@3954.6]
  wire [127:0] Z_70; // @[G128Multiplay.scala 38:7:@3953.4]
  wire  _T_1500; // @[G128Multiplay.scala 45:18:@3960.4]
  wire  _T_1502; // @[G128Multiplay.scala 45:22:@3961.4]
  wire [127:0] _T_1504; // @[G128Multiplay.scala 48:24:@3963.6]
  wire [127:0] _T_1508; // @[G128Multiplay.scala 51:31:@3969.6]
  wire [127:0] V_70; // @[G128Multiplay.scala 46:7:@3962.4]
  wire  _T_1510; // @[G128Multiplay.scala 37:16:@3973.4]
  wire [127:0] _T_1513; // @[G128Multiplay.scala 40:24:@3976.6]
  wire [127:0] Z_71; // @[G128Multiplay.scala 38:7:@3975.4]
  wire  _T_1514; // @[G128Multiplay.scala 45:18:@3982.4]
  wire  _T_1516; // @[G128Multiplay.scala 45:22:@3983.4]
  wire [127:0] _T_1518; // @[G128Multiplay.scala 48:24:@3985.6]
  wire [127:0] _T_1522; // @[G128Multiplay.scala 51:31:@3991.6]
  wire [127:0] V_71; // @[G128Multiplay.scala 46:7:@3984.4]
  wire  _T_1524; // @[G128Multiplay.scala 37:16:@3995.4]
  wire [127:0] _T_1527; // @[G128Multiplay.scala 40:24:@3998.6]
  wire [127:0] Z_72; // @[G128Multiplay.scala 38:7:@3997.4]
  wire  _T_1528; // @[G128Multiplay.scala 45:18:@4004.4]
  wire  _T_1530; // @[G128Multiplay.scala 45:22:@4005.4]
  wire [127:0] _T_1532; // @[G128Multiplay.scala 48:24:@4007.6]
  wire [127:0] _T_1536; // @[G128Multiplay.scala 51:31:@4013.6]
  wire [127:0] V_72; // @[G128Multiplay.scala 46:7:@4006.4]
  wire  _T_1538; // @[G128Multiplay.scala 37:16:@4017.4]
  wire [127:0] _T_1541; // @[G128Multiplay.scala 40:24:@4020.6]
  wire [127:0] Z_73; // @[G128Multiplay.scala 38:7:@4019.4]
  wire  _T_1542; // @[G128Multiplay.scala 45:18:@4026.4]
  wire  _T_1544; // @[G128Multiplay.scala 45:22:@4027.4]
  wire [127:0] _T_1546; // @[G128Multiplay.scala 48:24:@4029.6]
  wire [127:0] _T_1550; // @[G128Multiplay.scala 51:31:@4035.6]
  wire [127:0] V_73; // @[G128Multiplay.scala 46:7:@4028.4]
  wire  _T_1552; // @[G128Multiplay.scala 37:16:@4039.4]
  wire [127:0] _T_1555; // @[G128Multiplay.scala 40:24:@4042.6]
  wire [127:0] Z_74; // @[G128Multiplay.scala 38:7:@4041.4]
  wire  _T_1556; // @[G128Multiplay.scala 45:18:@4048.4]
  wire  _T_1558; // @[G128Multiplay.scala 45:22:@4049.4]
  wire [127:0] _T_1560; // @[G128Multiplay.scala 48:24:@4051.6]
  wire [127:0] _T_1564; // @[G128Multiplay.scala 51:31:@4057.6]
  wire [127:0] V_74; // @[G128Multiplay.scala 46:7:@4050.4]
  wire  _T_1566; // @[G128Multiplay.scala 37:16:@4061.4]
  wire [127:0] _T_1569; // @[G128Multiplay.scala 40:24:@4064.6]
  wire [127:0] Z_75; // @[G128Multiplay.scala 38:7:@4063.4]
  wire  _T_1570; // @[G128Multiplay.scala 45:18:@4070.4]
  wire  _T_1572; // @[G128Multiplay.scala 45:22:@4071.4]
  wire [127:0] _T_1574; // @[G128Multiplay.scala 48:24:@4073.6]
  wire [127:0] _T_1578; // @[G128Multiplay.scala 51:31:@4079.6]
  wire [127:0] V_75; // @[G128Multiplay.scala 46:7:@4072.4]
  wire  _T_1580; // @[G128Multiplay.scala 37:16:@4083.4]
  wire [127:0] _T_1583; // @[G128Multiplay.scala 40:24:@4086.6]
  wire [127:0] Z_76; // @[G128Multiplay.scala 38:7:@4085.4]
  wire  _T_1584; // @[G128Multiplay.scala 45:18:@4092.4]
  wire  _T_1586; // @[G128Multiplay.scala 45:22:@4093.4]
  wire [127:0] _T_1588; // @[G128Multiplay.scala 48:24:@4095.6]
  wire [127:0] _T_1592; // @[G128Multiplay.scala 51:31:@4101.6]
  wire [127:0] V_76; // @[G128Multiplay.scala 46:7:@4094.4]
  wire  _T_1594; // @[G128Multiplay.scala 37:16:@4105.4]
  wire [127:0] _T_1597; // @[G128Multiplay.scala 40:24:@4108.6]
  wire [127:0] Z_77; // @[G128Multiplay.scala 38:7:@4107.4]
  wire  _T_1598; // @[G128Multiplay.scala 45:18:@4114.4]
  wire  _T_1600; // @[G128Multiplay.scala 45:22:@4115.4]
  wire [127:0] _T_1602; // @[G128Multiplay.scala 48:24:@4117.6]
  wire [127:0] _T_1606; // @[G128Multiplay.scala 51:31:@4123.6]
  wire [127:0] V_77; // @[G128Multiplay.scala 46:7:@4116.4]
  wire  _T_1608; // @[G128Multiplay.scala 37:16:@4127.4]
  wire [127:0] _T_1611; // @[G128Multiplay.scala 40:24:@4130.6]
  wire [127:0] Z_78; // @[G128Multiplay.scala 38:7:@4129.4]
  wire  _T_1612; // @[G128Multiplay.scala 45:18:@4136.4]
  wire  _T_1614; // @[G128Multiplay.scala 45:22:@4137.4]
  wire [127:0] _T_1616; // @[G128Multiplay.scala 48:24:@4139.6]
  wire [127:0] _T_1620; // @[G128Multiplay.scala 51:31:@4145.6]
  wire [127:0] V_78; // @[G128Multiplay.scala 46:7:@4138.4]
  wire  _T_1622; // @[G128Multiplay.scala 37:16:@4149.4]
  wire [127:0] _T_1625; // @[G128Multiplay.scala 40:24:@4152.6]
  wire [127:0] Z_79; // @[G128Multiplay.scala 38:7:@4151.4]
  wire  _T_1626; // @[G128Multiplay.scala 45:18:@4158.4]
  wire  _T_1628; // @[G128Multiplay.scala 45:22:@4159.4]
  wire [127:0] _T_1630; // @[G128Multiplay.scala 48:24:@4161.6]
  wire [127:0] _T_1634; // @[G128Multiplay.scala 51:31:@4167.6]
  wire [127:0] V_79; // @[G128Multiplay.scala 46:7:@4160.4]
  wire  _T_1636; // @[G128Multiplay.scala 37:16:@4171.4]
  wire [127:0] _T_1639; // @[G128Multiplay.scala 40:24:@4174.6]
  wire [127:0] Z_80; // @[G128Multiplay.scala 38:7:@4173.4]
  wire  _T_1640; // @[G128Multiplay.scala 45:18:@4180.4]
  wire  _T_1642; // @[G128Multiplay.scala 45:22:@4181.4]
  wire [127:0] _T_1644; // @[G128Multiplay.scala 48:24:@4183.6]
  wire [127:0] _T_1648; // @[G128Multiplay.scala 51:31:@4189.6]
  wire [127:0] V_80; // @[G128Multiplay.scala 46:7:@4182.4]
  wire  _T_1650; // @[G128Multiplay.scala 37:16:@4193.4]
  wire [127:0] _T_1653; // @[G128Multiplay.scala 40:24:@4196.6]
  wire [127:0] Z_81; // @[G128Multiplay.scala 38:7:@4195.4]
  wire  _T_1654; // @[G128Multiplay.scala 45:18:@4202.4]
  wire  _T_1656; // @[G128Multiplay.scala 45:22:@4203.4]
  wire [127:0] _T_1658; // @[G128Multiplay.scala 48:24:@4205.6]
  wire [127:0] _T_1662; // @[G128Multiplay.scala 51:31:@4211.6]
  wire [127:0] V_81; // @[G128Multiplay.scala 46:7:@4204.4]
  wire  _T_1664; // @[G128Multiplay.scala 37:16:@4215.4]
  wire [127:0] _T_1667; // @[G128Multiplay.scala 40:24:@4218.6]
  wire [127:0] Z_82; // @[G128Multiplay.scala 38:7:@4217.4]
  wire  _T_1668; // @[G128Multiplay.scala 45:18:@4224.4]
  wire  _T_1670; // @[G128Multiplay.scala 45:22:@4225.4]
  wire [127:0] _T_1672; // @[G128Multiplay.scala 48:24:@4227.6]
  wire [127:0] _T_1676; // @[G128Multiplay.scala 51:31:@4233.6]
  wire [127:0] V_82; // @[G128Multiplay.scala 46:7:@4226.4]
  wire  _T_1678; // @[G128Multiplay.scala 37:16:@4237.4]
  wire [127:0] _T_1681; // @[G128Multiplay.scala 40:24:@4240.6]
  wire [127:0] Z_83; // @[G128Multiplay.scala 38:7:@4239.4]
  wire  _T_1682; // @[G128Multiplay.scala 45:18:@4246.4]
  wire  _T_1684; // @[G128Multiplay.scala 45:22:@4247.4]
  wire [127:0] _T_1686; // @[G128Multiplay.scala 48:24:@4249.6]
  wire [127:0] _T_1690; // @[G128Multiplay.scala 51:31:@4255.6]
  wire [127:0] V_83; // @[G128Multiplay.scala 46:7:@4248.4]
  wire  _T_1692; // @[G128Multiplay.scala 37:16:@4259.4]
  wire [127:0] _T_1695; // @[G128Multiplay.scala 40:24:@4262.6]
  wire [127:0] Z_84; // @[G128Multiplay.scala 38:7:@4261.4]
  wire  _T_1696; // @[G128Multiplay.scala 45:18:@4268.4]
  wire  _T_1698; // @[G128Multiplay.scala 45:22:@4269.4]
  wire [127:0] _T_1700; // @[G128Multiplay.scala 48:24:@4271.6]
  wire [127:0] _T_1704; // @[G128Multiplay.scala 51:31:@4277.6]
  wire [127:0] V_84; // @[G128Multiplay.scala 46:7:@4270.4]
  wire  _T_1706; // @[G128Multiplay.scala 37:16:@4281.4]
  wire [127:0] _T_1709; // @[G128Multiplay.scala 40:24:@4284.6]
  wire [127:0] Z_85; // @[G128Multiplay.scala 38:7:@4283.4]
  wire  _T_1710; // @[G128Multiplay.scala 45:18:@4290.4]
  wire  _T_1712; // @[G128Multiplay.scala 45:22:@4291.4]
  wire [127:0] _T_1714; // @[G128Multiplay.scala 48:24:@4293.6]
  wire [127:0] _T_1718; // @[G128Multiplay.scala 51:31:@4299.6]
  wire [127:0] V_85; // @[G128Multiplay.scala 46:7:@4292.4]
  wire  _T_1720; // @[G128Multiplay.scala 37:16:@4303.4]
  wire [127:0] _T_1723; // @[G128Multiplay.scala 40:24:@4306.6]
  wire [127:0] Z_86; // @[G128Multiplay.scala 38:7:@4305.4]
  wire  _T_1724; // @[G128Multiplay.scala 45:18:@4312.4]
  wire  _T_1726; // @[G128Multiplay.scala 45:22:@4313.4]
  wire [127:0] _T_1728; // @[G128Multiplay.scala 48:24:@4315.6]
  wire [127:0] _T_1732; // @[G128Multiplay.scala 51:31:@4321.6]
  wire [127:0] V_86; // @[G128Multiplay.scala 46:7:@4314.4]
  wire  _T_1734; // @[G128Multiplay.scala 37:16:@4325.4]
  wire [127:0] _T_1737; // @[G128Multiplay.scala 40:24:@4328.6]
  wire [127:0] Z_87; // @[G128Multiplay.scala 38:7:@4327.4]
  wire  _T_1738; // @[G128Multiplay.scala 45:18:@4334.4]
  wire  _T_1740; // @[G128Multiplay.scala 45:22:@4335.4]
  wire [127:0] _T_1742; // @[G128Multiplay.scala 48:24:@4337.6]
  wire [127:0] _T_1746; // @[G128Multiplay.scala 51:31:@4343.6]
  wire [127:0] V_87; // @[G128Multiplay.scala 46:7:@4336.4]
  wire  _T_1748; // @[G128Multiplay.scala 37:16:@4347.4]
  wire [127:0] _T_1751; // @[G128Multiplay.scala 40:24:@4350.6]
  wire [127:0] Z_88; // @[G128Multiplay.scala 38:7:@4349.4]
  wire  _T_1752; // @[G128Multiplay.scala 45:18:@4356.4]
  wire  _T_1754; // @[G128Multiplay.scala 45:22:@4357.4]
  wire [127:0] _T_1756; // @[G128Multiplay.scala 48:24:@4359.6]
  wire [127:0] _T_1760; // @[G128Multiplay.scala 51:31:@4365.6]
  wire [127:0] V_88; // @[G128Multiplay.scala 46:7:@4358.4]
  wire  _T_1762; // @[G128Multiplay.scala 37:16:@4369.4]
  wire [127:0] _T_1765; // @[G128Multiplay.scala 40:24:@4372.6]
  wire [127:0] Z_89; // @[G128Multiplay.scala 38:7:@4371.4]
  wire  _T_1766; // @[G128Multiplay.scala 45:18:@4378.4]
  wire  _T_1768; // @[G128Multiplay.scala 45:22:@4379.4]
  wire [127:0] _T_1770; // @[G128Multiplay.scala 48:24:@4381.6]
  wire [127:0] _T_1774; // @[G128Multiplay.scala 51:31:@4387.6]
  wire [127:0] V_89; // @[G128Multiplay.scala 46:7:@4380.4]
  wire  _T_1776; // @[G128Multiplay.scala 37:16:@4391.4]
  wire [127:0] _T_1779; // @[G128Multiplay.scala 40:24:@4394.6]
  wire [127:0] Z_90; // @[G128Multiplay.scala 38:7:@4393.4]
  wire  _T_1780; // @[G128Multiplay.scala 45:18:@4400.4]
  wire  _T_1782; // @[G128Multiplay.scala 45:22:@4401.4]
  wire [127:0] _T_1784; // @[G128Multiplay.scala 48:24:@4403.6]
  wire [127:0] _T_1788; // @[G128Multiplay.scala 51:31:@4409.6]
  wire [127:0] V_90; // @[G128Multiplay.scala 46:7:@4402.4]
  wire  _T_1790; // @[G128Multiplay.scala 37:16:@4413.4]
  wire [127:0] _T_1793; // @[G128Multiplay.scala 40:24:@4416.6]
  wire [127:0] Z_91; // @[G128Multiplay.scala 38:7:@4415.4]
  wire  _T_1794; // @[G128Multiplay.scala 45:18:@4422.4]
  wire  _T_1796; // @[G128Multiplay.scala 45:22:@4423.4]
  wire [127:0] _T_1798; // @[G128Multiplay.scala 48:24:@4425.6]
  wire [127:0] _T_1802; // @[G128Multiplay.scala 51:31:@4431.6]
  wire [127:0] V_91; // @[G128Multiplay.scala 46:7:@4424.4]
  wire  _T_1804; // @[G128Multiplay.scala 37:16:@4435.4]
  wire [127:0] _T_1807; // @[G128Multiplay.scala 40:24:@4438.6]
  wire [127:0] Z_92; // @[G128Multiplay.scala 38:7:@4437.4]
  wire  _T_1808; // @[G128Multiplay.scala 45:18:@4444.4]
  wire  _T_1810; // @[G128Multiplay.scala 45:22:@4445.4]
  wire [127:0] _T_1812; // @[G128Multiplay.scala 48:24:@4447.6]
  wire [127:0] _T_1816; // @[G128Multiplay.scala 51:31:@4453.6]
  wire [127:0] V_92; // @[G128Multiplay.scala 46:7:@4446.4]
  wire  _T_1818; // @[G128Multiplay.scala 37:16:@4457.4]
  wire [127:0] _T_1821; // @[G128Multiplay.scala 40:24:@4460.6]
  wire [127:0] Z_93; // @[G128Multiplay.scala 38:7:@4459.4]
  wire  _T_1822; // @[G128Multiplay.scala 45:18:@4466.4]
  wire  _T_1824; // @[G128Multiplay.scala 45:22:@4467.4]
  wire [127:0] _T_1826; // @[G128Multiplay.scala 48:24:@4469.6]
  wire [127:0] _T_1830; // @[G128Multiplay.scala 51:31:@4475.6]
  wire [127:0] V_93; // @[G128Multiplay.scala 46:7:@4468.4]
  wire  _T_1832; // @[G128Multiplay.scala 37:16:@4479.4]
  wire [127:0] _T_1835; // @[G128Multiplay.scala 40:24:@4482.6]
  wire [127:0] Z_94; // @[G128Multiplay.scala 38:7:@4481.4]
  wire  _T_1836; // @[G128Multiplay.scala 45:18:@4488.4]
  wire  _T_1838; // @[G128Multiplay.scala 45:22:@4489.4]
  wire [127:0] _T_1840; // @[G128Multiplay.scala 48:24:@4491.6]
  wire [127:0] _T_1844; // @[G128Multiplay.scala 51:31:@4497.6]
  wire [127:0] V_94; // @[G128Multiplay.scala 46:7:@4490.4]
  wire  _T_1846; // @[G128Multiplay.scala 37:16:@4501.4]
  wire [127:0] _T_1849; // @[G128Multiplay.scala 40:24:@4504.6]
  wire [127:0] Z_95; // @[G128Multiplay.scala 38:7:@4503.4]
  wire  _T_1850; // @[G128Multiplay.scala 45:18:@4510.4]
  wire  _T_1852; // @[G128Multiplay.scala 45:22:@4511.4]
  wire [127:0] _T_1854; // @[G128Multiplay.scala 48:24:@4513.6]
  wire [127:0] _T_1858; // @[G128Multiplay.scala 51:31:@4519.6]
  wire [127:0] V_95; // @[G128Multiplay.scala 46:7:@4512.4]
  wire  _T_1860; // @[G128Multiplay.scala 37:16:@4523.4]
  wire [127:0] _T_1863; // @[G128Multiplay.scala 40:24:@4526.6]
  wire [127:0] Z_96; // @[G128Multiplay.scala 38:7:@4525.4]
  wire  _T_1864; // @[G128Multiplay.scala 45:18:@4532.4]
  wire  _T_1866; // @[G128Multiplay.scala 45:22:@4533.4]
  wire [127:0] _T_1868; // @[G128Multiplay.scala 48:24:@4535.6]
  wire [127:0] _T_1872; // @[G128Multiplay.scala 51:31:@4541.6]
  wire [127:0] V_96; // @[G128Multiplay.scala 46:7:@4534.4]
  wire  _T_1874; // @[G128Multiplay.scala 37:16:@4545.4]
  wire [127:0] _T_1877; // @[G128Multiplay.scala 40:24:@4548.6]
  wire [127:0] Z_97; // @[G128Multiplay.scala 38:7:@4547.4]
  wire  _T_1878; // @[G128Multiplay.scala 45:18:@4554.4]
  wire  _T_1880; // @[G128Multiplay.scala 45:22:@4555.4]
  wire [127:0] _T_1882; // @[G128Multiplay.scala 48:24:@4557.6]
  wire [127:0] _T_1886; // @[G128Multiplay.scala 51:31:@4563.6]
  wire [127:0] V_97; // @[G128Multiplay.scala 46:7:@4556.4]
  wire  _T_1888; // @[G128Multiplay.scala 37:16:@4567.4]
  wire [127:0] _T_1891; // @[G128Multiplay.scala 40:24:@4570.6]
  wire [127:0] Z_98; // @[G128Multiplay.scala 38:7:@4569.4]
  wire  _T_1892; // @[G128Multiplay.scala 45:18:@4576.4]
  wire  _T_1894; // @[G128Multiplay.scala 45:22:@4577.4]
  wire [127:0] _T_1896; // @[G128Multiplay.scala 48:24:@4579.6]
  wire [127:0] _T_1900; // @[G128Multiplay.scala 51:31:@4585.6]
  wire [127:0] V_98; // @[G128Multiplay.scala 46:7:@4578.4]
  wire  _T_1902; // @[G128Multiplay.scala 37:16:@4589.4]
  wire [127:0] _T_1905; // @[G128Multiplay.scala 40:24:@4592.6]
  wire [127:0] Z_99; // @[G128Multiplay.scala 38:7:@4591.4]
  wire  _T_1906; // @[G128Multiplay.scala 45:18:@4598.4]
  wire  _T_1908; // @[G128Multiplay.scala 45:22:@4599.4]
  wire [127:0] _T_1910; // @[G128Multiplay.scala 48:24:@4601.6]
  wire [127:0] _T_1914; // @[G128Multiplay.scala 51:31:@4607.6]
  wire [127:0] V_99; // @[G128Multiplay.scala 46:7:@4600.4]
  wire  _T_1916; // @[G128Multiplay.scala 37:16:@4611.4]
  wire [127:0] _T_1919; // @[G128Multiplay.scala 40:24:@4614.6]
  wire [127:0] Z_100; // @[G128Multiplay.scala 38:7:@4613.4]
  wire  _T_1920; // @[G128Multiplay.scala 45:18:@4620.4]
  wire  _T_1922; // @[G128Multiplay.scala 45:22:@4621.4]
  wire [127:0] _T_1924; // @[G128Multiplay.scala 48:24:@4623.6]
  wire [127:0] _T_1928; // @[G128Multiplay.scala 51:31:@4629.6]
  wire [127:0] V_100; // @[G128Multiplay.scala 46:7:@4622.4]
  wire  _T_1930; // @[G128Multiplay.scala 37:16:@4633.4]
  wire [127:0] _T_1933; // @[G128Multiplay.scala 40:24:@4636.6]
  wire [127:0] Z_101; // @[G128Multiplay.scala 38:7:@4635.4]
  wire  _T_1934; // @[G128Multiplay.scala 45:18:@4642.4]
  wire  _T_1936; // @[G128Multiplay.scala 45:22:@4643.4]
  wire [127:0] _T_1938; // @[G128Multiplay.scala 48:24:@4645.6]
  wire [127:0] _T_1942; // @[G128Multiplay.scala 51:31:@4651.6]
  wire [127:0] V_101; // @[G128Multiplay.scala 46:7:@4644.4]
  wire  _T_1944; // @[G128Multiplay.scala 37:16:@4655.4]
  wire [127:0] _T_1947; // @[G128Multiplay.scala 40:24:@4658.6]
  wire [127:0] Z_102; // @[G128Multiplay.scala 38:7:@4657.4]
  wire  _T_1948; // @[G128Multiplay.scala 45:18:@4664.4]
  wire  _T_1950; // @[G128Multiplay.scala 45:22:@4665.4]
  wire [127:0] _T_1952; // @[G128Multiplay.scala 48:24:@4667.6]
  wire [127:0] _T_1956; // @[G128Multiplay.scala 51:31:@4673.6]
  wire [127:0] V_102; // @[G128Multiplay.scala 46:7:@4666.4]
  wire  _T_1958; // @[G128Multiplay.scala 37:16:@4677.4]
  wire [127:0] _T_1961; // @[G128Multiplay.scala 40:24:@4680.6]
  wire [127:0] Z_103; // @[G128Multiplay.scala 38:7:@4679.4]
  wire  _T_1962; // @[G128Multiplay.scala 45:18:@4686.4]
  wire  _T_1964; // @[G128Multiplay.scala 45:22:@4687.4]
  wire [127:0] _T_1966; // @[G128Multiplay.scala 48:24:@4689.6]
  wire [127:0] _T_1970; // @[G128Multiplay.scala 51:31:@4695.6]
  wire [127:0] V_103; // @[G128Multiplay.scala 46:7:@4688.4]
  wire  _T_1972; // @[G128Multiplay.scala 37:16:@4699.4]
  wire [127:0] _T_1975; // @[G128Multiplay.scala 40:24:@4702.6]
  wire [127:0] Z_104; // @[G128Multiplay.scala 38:7:@4701.4]
  wire  _T_1976; // @[G128Multiplay.scala 45:18:@4708.4]
  wire  _T_1978; // @[G128Multiplay.scala 45:22:@4709.4]
  wire [127:0] _T_1980; // @[G128Multiplay.scala 48:24:@4711.6]
  wire [127:0] _T_1984; // @[G128Multiplay.scala 51:31:@4717.6]
  wire [127:0] V_104; // @[G128Multiplay.scala 46:7:@4710.4]
  wire  _T_1986; // @[G128Multiplay.scala 37:16:@4721.4]
  wire [127:0] _T_1989; // @[G128Multiplay.scala 40:24:@4724.6]
  wire [127:0] Z_105; // @[G128Multiplay.scala 38:7:@4723.4]
  wire  _T_1990; // @[G128Multiplay.scala 45:18:@4730.4]
  wire  _T_1992; // @[G128Multiplay.scala 45:22:@4731.4]
  wire [127:0] _T_1994; // @[G128Multiplay.scala 48:24:@4733.6]
  wire [127:0] _T_1998; // @[G128Multiplay.scala 51:31:@4739.6]
  wire [127:0] V_105; // @[G128Multiplay.scala 46:7:@4732.4]
  wire  _T_2000; // @[G128Multiplay.scala 37:16:@4743.4]
  wire [127:0] _T_2003; // @[G128Multiplay.scala 40:24:@4746.6]
  wire [127:0] Z_106; // @[G128Multiplay.scala 38:7:@4745.4]
  wire  _T_2004; // @[G128Multiplay.scala 45:18:@4752.4]
  wire  _T_2006; // @[G128Multiplay.scala 45:22:@4753.4]
  wire [127:0] _T_2008; // @[G128Multiplay.scala 48:24:@4755.6]
  wire [127:0] _T_2012; // @[G128Multiplay.scala 51:31:@4761.6]
  wire [127:0] V_106; // @[G128Multiplay.scala 46:7:@4754.4]
  wire  _T_2014; // @[G128Multiplay.scala 37:16:@4765.4]
  wire [127:0] _T_2017; // @[G128Multiplay.scala 40:24:@4768.6]
  wire [127:0] Z_107; // @[G128Multiplay.scala 38:7:@4767.4]
  wire  _T_2018; // @[G128Multiplay.scala 45:18:@4774.4]
  wire  _T_2020; // @[G128Multiplay.scala 45:22:@4775.4]
  wire [127:0] _T_2022; // @[G128Multiplay.scala 48:24:@4777.6]
  wire [127:0] _T_2026; // @[G128Multiplay.scala 51:31:@4783.6]
  wire [127:0] V_107; // @[G128Multiplay.scala 46:7:@4776.4]
  wire  _T_2028; // @[G128Multiplay.scala 37:16:@4787.4]
  wire [127:0] _T_2031; // @[G128Multiplay.scala 40:24:@4790.6]
  wire [127:0] Z_108; // @[G128Multiplay.scala 38:7:@4789.4]
  wire  _T_2032; // @[G128Multiplay.scala 45:18:@4796.4]
  wire  _T_2034; // @[G128Multiplay.scala 45:22:@4797.4]
  wire [127:0] _T_2036; // @[G128Multiplay.scala 48:24:@4799.6]
  wire [127:0] _T_2040; // @[G128Multiplay.scala 51:31:@4805.6]
  wire [127:0] V_108; // @[G128Multiplay.scala 46:7:@4798.4]
  wire  _T_2042; // @[G128Multiplay.scala 37:16:@4809.4]
  wire [127:0] _T_2045; // @[G128Multiplay.scala 40:24:@4812.6]
  wire [127:0] Z_109; // @[G128Multiplay.scala 38:7:@4811.4]
  wire  _T_2046; // @[G128Multiplay.scala 45:18:@4818.4]
  wire  _T_2048; // @[G128Multiplay.scala 45:22:@4819.4]
  wire [127:0] _T_2050; // @[G128Multiplay.scala 48:24:@4821.6]
  wire [127:0] _T_2054; // @[G128Multiplay.scala 51:31:@4827.6]
  wire [127:0] V_109; // @[G128Multiplay.scala 46:7:@4820.4]
  wire  _T_2056; // @[G128Multiplay.scala 37:16:@4831.4]
  wire [127:0] _T_2059; // @[G128Multiplay.scala 40:24:@4834.6]
  wire [127:0] Z_110; // @[G128Multiplay.scala 38:7:@4833.4]
  wire  _T_2060; // @[G128Multiplay.scala 45:18:@4840.4]
  wire  _T_2062; // @[G128Multiplay.scala 45:22:@4841.4]
  wire [127:0] _T_2064; // @[G128Multiplay.scala 48:24:@4843.6]
  wire [127:0] _T_2068; // @[G128Multiplay.scala 51:31:@4849.6]
  wire [127:0] V_110; // @[G128Multiplay.scala 46:7:@4842.4]
  wire  _T_2070; // @[G128Multiplay.scala 37:16:@4853.4]
  wire [127:0] _T_2073; // @[G128Multiplay.scala 40:24:@4856.6]
  wire [127:0] Z_111; // @[G128Multiplay.scala 38:7:@4855.4]
  wire  _T_2074; // @[G128Multiplay.scala 45:18:@4862.4]
  wire  _T_2076; // @[G128Multiplay.scala 45:22:@4863.4]
  wire [127:0] _T_2078; // @[G128Multiplay.scala 48:24:@4865.6]
  wire [127:0] _T_2082; // @[G128Multiplay.scala 51:31:@4871.6]
  wire [127:0] V_111; // @[G128Multiplay.scala 46:7:@4864.4]
  wire  _T_2084; // @[G128Multiplay.scala 37:16:@4875.4]
  wire [127:0] _T_2087; // @[G128Multiplay.scala 40:24:@4878.6]
  wire [127:0] Z_112; // @[G128Multiplay.scala 38:7:@4877.4]
  wire  _T_2088; // @[G128Multiplay.scala 45:18:@4884.4]
  wire  _T_2090; // @[G128Multiplay.scala 45:22:@4885.4]
  wire [127:0] _T_2092; // @[G128Multiplay.scala 48:24:@4887.6]
  wire [127:0] _T_2096; // @[G128Multiplay.scala 51:31:@4893.6]
  wire [127:0] V_112; // @[G128Multiplay.scala 46:7:@4886.4]
  wire  _T_2098; // @[G128Multiplay.scala 37:16:@4897.4]
  wire [127:0] _T_2101; // @[G128Multiplay.scala 40:24:@4900.6]
  wire [127:0] Z_113; // @[G128Multiplay.scala 38:7:@4899.4]
  wire  _T_2102; // @[G128Multiplay.scala 45:18:@4906.4]
  wire  _T_2104; // @[G128Multiplay.scala 45:22:@4907.4]
  wire [127:0] _T_2106; // @[G128Multiplay.scala 48:24:@4909.6]
  wire [127:0] _T_2110; // @[G128Multiplay.scala 51:31:@4915.6]
  wire [127:0] V_113; // @[G128Multiplay.scala 46:7:@4908.4]
  wire  _T_2112; // @[G128Multiplay.scala 37:16:@4919.4]
  wire [127:0] _T_2115; // @[G128Multiplay.scala 40:24:@4922.6]
  wire [127:0] Z_114; // @[G128Multiplay.scala 38:7:@4921.4]
  wire  _T_2116; // @[G128Multiplay.scala 45:18:@4928.4]
  wire  _T_2118; // @[G128Multiplay.scala 45:22:@4929.4]
  wire [127:0] _T_2120; // @[G128Multiplay.scala 48:24:@4931.6]
  wire [127:0] _T_2124; // @[G128Multiplay.scala 51:31:@4937.6]
  wire [127:0] V_114; // @[G128Multiplay.scala 46:7:@4930.4]
  wire  _T_2126; // @[G128Multiplay.scala 37:16:@4941.4]
  wire [127:0] _T_2129; // @[G128Multiplay.scala 40:24:@4944.6]
  wire [127:0] Z_115; // @[G128Multiplay.scala 38:7:@4943.4]
  wire  _T_2130; // @[G128Multiplay.scala 45:18:@4950.4]
  wire  _T_2132; // @[G128Multiplay.scala 45:22:@4951.4]
  wire [127:0] _T_2134; // @[G128Multiplay.scala 48:24:@4953.6]
  wire [127:0] _T_2138; // @[G128Multiplay.scala 51:31:@4959.6]
  wire [127:0] V_115; // @[G128Multiplay.scala 46:7:@4952.4]
  wire  _T_2140; // @[G128Multiplay.scala 37:16:@4963.4]
  wire [127:0] _T_2143; // @[G128Multiplay.scala 40:24:@4966.6]
  wire [127:0] Z_116; // @[G128Multiplay.scala 38:7:@4965.4]
  wire  _T_2144; // @[G128Multiplay.scala 45:18:@4972.4]
  wire  _T_2146; // @[G128Multiplay.scala 45:22:@4973.4]
  wire [127:0] _T_2148; // @[G128Multiplay.scala 48:24:@4975.6]
  wire [127:0] _T_2152; // @[G128Multiplay.scala 51:31:@4981.6]
  wire [127:0] V_116; // @[G128Multiplay.scala 46:7:@4974.4]
  wire  _T_2154; // @[G128Multiplay.scala 37:16:@4985.4]
  wire [127:0] _T_2157; // @[G128Multiplay.scala 40:24:@4988.6]
  wire [127:0] Z_117; // @[G128Multiplay.scala 38:7:@4987.4]
  wire  _T_2158; // @[G128Multiplay.scala 45:18:@4994.4]
  wire  _T_2160; // @[G128Multiplay.scala 45:22:@4995.4]
  wire [127:0] _T_2162; // @[G128Multiplay.scala 48:24:@4997.6]
  wire [127:0] _T_2166; // @[G128Multiplay.scala 51:31:@5003.6]
  wire [127:0] V_117; // @[G128Multiplay.scala 46:7:@4996.4]
  wire  _T_2168; // @[G128Multiplay.scala 37:16:@5007.4]
  wire [127:0] _T_2171; // @[G128Multiplay.scala 40:24:@5010.6]
  wire [127:0] Z_118; // @[G128Multiplay.scala 38:7:@5009.4]
  wire  _T_2172; // @[G128Multiplay.scala 45:18:@5016.4]
  wire  _T_2174; // @[G128Multiplay.scala 45:22:@5017.4]
  wire [127:0] _T_2176; // @[G128Multiplay.scala 48:24:@5019.6]
  wire [127:0] _T_2180; // @[G128Multiplay.scala 51:31:@5025.6]
  wire [127:0] V_118; // @[G128Multiplay.scala 46:7:@5018.4]
  wire  _T_2182; // @[G128Multiplay.scala 37:16:@5029.4]
  wire [127:0] _T_2185; // @[G128Multiplay.scala 40:24:@5032.6]
  wire [127:0] Z_119; // @[G128Multiplay.scala 38:7:@5031.4]
  wire  _T_2186; // @[G128Multiplay.scala 45:18:@5038.4]
  wire  _T_2188; // @[G128Multiplay.scala 45:22:@5039.4]
  wire [127:0] _T_2190; // @[G128Multiplay.scala 48:24:@5041.6]
  wire [127:0] _T_2194; // @[G128Multiplay.scala 51:31:@5047.6]
  wire [127:0] V_119; // @[G128Multiplay.scala 46:7:@5040.4]
  wire  _T_2196; // @[G128Multiplay.scala 37:16:@5051.4]
  wire [127:0] _T_2199; // @[G128Multiplay.scala 40:24:@5054.6]
  wire [127:0] Z_120; // @[G128Multiplay.scala 38:7:@5053.4]
  wire  _T_2200; // @[G128Multiplay.scala 45:18:@5060.4]
  wire  _T_2202; // @[G128Multiplay.scala 45:22:@5061.4]
  wire [127:0] _T_2204; // @[G128Multiplay.scala 48:24:@5063.6]
  wire [127:0] _T_2208; // @[G128Multiplay.scala 51:31:@5069.6]
  wire [127:0] V_120; // @[G128Multiplay.scala 46:7:@5062.4]
  wire  _T_2210; // @[G128Multiplay.scala 37:16:@5073.4]
  wire [127:0] _T_2213; // @[G128Multiplay.scala 40:24:@5076.6]
  wire [127:0] Z_121; // @[G128Multiplay.scala 38:7:@5075.4]
  wire  _T_2214; // @[G128Multiplay.scala 45:18:@5082.4]
  wire  _T_2216; // @[G128Multiplay.scala 45:22:@5083.4]
  wire [127:0] _T_2218; // @[G128Multiplay.scala 48:24:@5085.6]
  wire [127:0] _T_2222; // @[G128Multiplay.scala 51:31:@5091.6]
  wire [127:0] V_121; // @[G128Multiplay.scala 46:7:@5084.4]
  wire  _T_2224; // @[G128Multiplay.scala 37:16:@5095.4]
  wire [127:0] _T_2227; // @[G128Multiplay.scala 40:24:@5098.6]
  wire [127:0] Z_122; // @[G128Multiplay.scala 38:7:@5097.4]
  wire  _T_2228; // @[G128Multiplay.scala 45:18:@5104.4]
  wire  _T_2230; // @[G128Multiplay.scala 45:22:@5105.4]
  wire [127:0] _T_2232; // @[G128Multiplay.scala 48:24:@5107.6]
  wire [127:0] _T_2236; // @[G128Multiplay.scala 51:31:@5113.6]
  wire [127:0] V_122; // @[G128Multiplay.scala 46:7:@5106.4]
  wire  _T_2238; // @[G128Multiplay.scala 37:16:@5117.4]
  wire [127:0] _T_2241; // @[G128Multiplay.scala 40:24:@5120.6]
  wire [127:0] Z_123; // @[G128Multiplay.scala 38:7:@5119.4]
  wire  _T_2242; // @[G128Multiplay.scala 45:18:@5126.4]
  wire  _T_2244; // @[G128Multiplay.scala 45:22:@5127.4]
  wire [127:0] _T_2246; // @[G128Multiplay.scala 48:24:@5129.6]
  wire [127:0] _T_2250; // @[G128Multiplay.scala 51:31:@5135.6]
  wire [127:0] V_123; // @[G128Multiplay.scala 46:7:@5128.4]
  wire  _T_2252; // @[G128Multiplay.scala 37:16:@5139.4]
  wire [127:0] _T_2255; // @[G128Multiplay.scala 40:24:@5142.6]
  wire [127:0] Z_124; // @[G128Multiplay.scala 38:7:@5141.4]
  wire  _T_2256; // @[G128Multiplay.scala 45:18:@5148.4]
  wire  _T_2258; // @[G128Multiplay.scala 45:22:@5149.4]
  wire [127:0] _T_2260; // @[G128Multiplay.scala 48:24:@5151.6]
  wire [127:0] _T_2264; // @[G128Multiplay.scala 51:31:@5157.6]
  wire [127:0] V_124; // @[G128Multiplay.scala 46:7:@5150.4]
  wire  _T_2266; // @[G128Multiplay.scala 37:16:@5161.4]
  wire [127:0] _T_2269; // @[G128Multiplay.scala 40:24:@5164.6]
  wire [127:0] Z_125; // @[G128Multiplay.scala 38:7:@5163.4]
  wire  _T_2270; // @[G128Multiplay.scala 45:18:@5170.4]
  wire  _T_2272; // @[G128Multiplay.scala 45:22:@5171.4]
  wire [127:0] _T_2274; // @[G128Multiplay.scala 48:24:@5173.6]
  wire [127:0] _T_2278; // @[G128Multiplay.scala 51:31:@5179.6]
  wire [127:0] V_125; // @[G128Multiplay.scala 46:7:@5172.4]
  wire  _T_2280; // @[G128Multiplay.scala 37:16:@5183.4]
  wire [127:0] _T_2283; // @[G128Multiplay.scala 40:24:@5186.6]
  wire [127:0] Z_126; // @[G128Multiplay.scala 38:7:@5185.4]
  wire  _T_2284; // @[G128Multiplay.scala 45:18:@5192.4]
  wire  _T_2286; // @[G128Multiplay.scala 45:22:@5193.4]
  wire [127:0] _T_2288; // @[G128Multiplay.scala 48:24:@5195.6]
  wire [127:0] _T_2292; // @[G128Multiplay.scala 51:31:@5201.6]
  wire [127:0] V_126; // @[G128Multiplay.scala 46:7:@5194.4]
  wire  _T_2294; // @[G128Multiplay.scala 37:16:@5205.4]
  wire [127:0] _T_2297; // @[G128Multiplay.scala 40:24:@5208.6]
  wire [127:0] Z_127; // @[G128Multiplay.scala 38:7:@5207.4]
  wire  _T_2298; // @[G128Multiplay.scala 45:18:@5214.4]
  wire  _T_2300; // @[G128Multiplay.scala 45:22:@5215.4]
  wire [127:0] _T_2302; // @[G128Multiplay.scala 48:24:@5217.6]
  wire [127:0] _T_2306; // @[G128Multiplay.scala 51:31:@5223.6]
  wire [127:0] V_127; // @[G128Multiplay.scala 46:7:@5216.4]
  wire  _T_2308; // @[G128Multiplay.scala 37:16:@5227.4]
  wire [127:0] _T_2311; // @[G128Multiplay.scala 40:24:@5230.6]
  wire [127:0] Z_128; // @[G128Multiplay.scala 38:7:@5229.4]
  assign _T_530 = io_y[127]; // @[G128Multiplay.scala 37:16:@2433.4]
  assign Z_1 = _T_530 ? io_x : 128'h0; // @[G128Multiplay.scala 38:7:@2435.4]
  assign _T_534 = io_x[0]; // @[G128Multiplay.scala 45:18:@2442.4]
  assign _T_536 = _T_534 == 1'h0; // @[G128Multiplay.scala 45:22:@2443.4]
  assign _T_538 = io_x >> 1'h1; // @[G128Multiplay.scala 48:24:@2445.6]
  assign _T_542 = _T_538 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2451.6]
  assign V_1 = _T_536 ? _T_538 : _T_542; // @[G128Multiplay.scala 46:7:@2444.4]
  assign _T_544 = io_y[126]; // @[G128Multiplay.scala 37:16:@2455.4]
  assign _T_547 = Z_1 ^ V_1; // @[G128Multiplay.scala 40:24:@2458.6]
  assign Z_2 = _T_544 ? _T_547 : Z_1; // @[G128Multiplay.scala 38:7:@2457.4]
  assign _T_548 = V_1[0]; // @[G128Multiplay.scala 45:18:@2464.4]
  assign _T_550 = _T_548 == 1'h0; // @[G128Multiplay.scala 45:22:@2465.4]
  assign _T_552 = V_1 >> 1'h1; // @[G128Multiplay.scala 48:24:@2467.6]
  assign _T_556 = _T_552 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2473.6]
  assign V_2 = _T_550 ? _T_552 : _T_556; // @[G128Multiplay.scala 46:7:@2466.4]
  assign _T_558 = io_y[125]; // @[G128Multiplay.scala 37:16:@2477.4]
  assign _T_561 = Z_2 ^ V_2; // @[G128Multiplay.scala 40:24:@2480.6]
  assign Z_3 = _T_558 ? _T_561 : Z_2; // @[G128Multiplay.scala 38:7:@2479.4]
  assign _T_562 = V_2[0]; // @[G128Multiplay.scala 45:18:@2486.4]
  assign _T_564 = _T_562 == 1'h0; // @[G128Multiplay.scala 45:22:@2487.4]
  assign _T_566 = V_2 >> 1'h1; // @[G128Multiplay.scala 48:24:@2489.6]
  assign _T_570 = _T_566 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2495.6]
  assign V_3 = _T_564 ? _T_566 : _T_570; // @[G128Multiplay.scala 46:7:@2488.4]
  assign _T_572 = io_y[124]; // @[G128Multiplay.scala 37:16:@2499.4]
  assign _T_575 = Z_3 ^ V_3; // @[G128Multiplay.scala 40:24:@2502.6]
  assign Z_4 = _T_572 ? _T_575 : Z_3; // @[G128Multiplay.scala 38:7:@2501.4]
  assign _T_576 = V_3[0]; // @[G128Multiplay.scala 45:18:@2508.4]
  assign _T_578 = _T_576 == 1'h0; // @[G128Multiplay.scala 45:22:@2509.4]
  assign _T_580 = V_3 >> 1'h1; // @[G128Multiplay.scala 48:24:@2511.6]
  assign _T_584 = _T_580 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2517.6]
  assign V_4 = _T_578 ? _T_580 : _T_584; // @[G128Multiplay.scala 46:7:@2510.4]
  assign _T_586 = io_y[123]; // @[G128Multiplay.scala 37:16:@2521.4]
  assign _T_589 = Z_4 ^ V_4; // @[G128Multiplay.scala 40:24:@2524.6]
  assign Z_5 = _T_586 ? _T_589 : Z_4; // @[G128Multiplay.scala 38:7:@2523.4]
  assign _T_590 = V_4[0]; // @[G128Multiplay.scala 45:18:@2530.4]
  assign _T_592 = _T_590 == 1'h0; // @[G128Multiplay.scala 45:22:@2531.4]
  assign _T_594 = V_4 >> 1'h1; // @[G128Multiplay.scala 48:24:@2533.6]
  assign _T_598 = _T_594 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2539.6]
  assign V_5 = _T_592 ? _T_594 : _T_598; // @[G128Multiplay.scala 46:7:@2532.4]
  assign _T_600 = io_y[122]; // @[G128Multiplay.scala 37:16:@2543.4]
  assign _T_603 = Z_5 ^ V_5; // @[G128Multiplay.scala 40:24:@2546.6]
  assign Z_6 = _T_600 ? _T_603 : Z_5; // @[G128Multiplay.scala 38:7:@2545.4]
  assign _T_604 = V_5[0]; // @[G128Multiplay.scala 45:18:@2552.4]
  assign _T_606 = _T_604 == 1'h0; // @[G128Multiplay.scala 45:22:@2553.4]
  assign _T_608 = V_5 >> 1'h1; // @[G128Multiplay.scala 48:24:@2555.6]
  assign _T_612 = _T_608 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2561.6]
  assign V_6 = _T_606 ? _T_608 : _T_612; // @[G128Multiplay.scala 46:7:@2554.4]
  assign _T_614 = io_y[121]; // @[G128Multiplay.scala 37:16:@2565.4]
  assign _T_617 = Z_6 ^ V_6; // @[G128Multiplay.scala 40:24:@2568.6]
  assign Z_7 = _T_614 ? _T_617 : Z_6; // @[G128Multiplay.scala 38:7:@2567.4]
  assign _T_618 = V_6[0]; // @[G128Multiplay.scala 45:18:@2574.4]
  assign _T_620 = _T_618 == 1'h0; // @[G128Multiplay.scala 45:22:@2575.4]
  assign _T_622 = V_6 >> 1'h1; // @[G128Multiplay.scala 48:24:@2577.6]
  assign _T_626 = _T_622 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2583.6]
  assign V_7 = _T_620 ? _T_622 : _T_626; // @[G128Multiplay.scala 46:7:@2576.4]
  assign _T_628 = io_y[120]; // @[G128Multiplay.scala 37:16:@2587.4]
  assign _T_631 = Z_7 ^ V_7; // @[G128Multiplay.scala 40:24:@2590.6]
  assign Z_8 = _T_628 ? _T_631 : Z_7; // @[G128Multiplay.scala 38:7:@2589.4]
  assign _T_632 = V_7[0]; // @[G128Multiplay.scala 45:18:@2596.4]
  assign _T_634 = _T_632 == 1'h0; // @[G128Multiplay.scala 45:22:@2597.4]
  assign _T_636 = V_7 >> 1'h1; // @[G128Multiplay.scala 48:24:@2599.6]
  assign _T_640 = _T_636 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2605.6]
  assign V_8 = _T_634 ? _T_636 : _T_640; // @[G128Multiplay.scala 46:7:@2598.4]
  assign _T_642 = io_y[119]; // @[G128Multiplay.scala 37:16:@2609.4]
  assign _T_645 = Z_8 ^ V_8; // @[G128Multiplay.scala 40:24:@2612.6]
  assign Z_9 = _T_642 ? _T_645 : Z_8; // @[G128Multiplay.scala 38:7:@2611.4]
  assign _T_646 = V_8[0]; // @[G128Multiplay.scala 45:18:@2618.4]
  assign _T_648 = _T_646 == 1'h0; // @[G128Multiplay.scala 45:22:@2619.4]
  assign _T_650 = V_8 >> 1'h1; // @[G128Multiplay.scala 48:24:@2621.6]
  assign _T_654 = _T_650 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2627.6]
  assign V_9 = _T_648 ? _T_650 : _T_654; // @[G128Multiplay.scala 46:7:@2620.4]
  assign _T_656 = io_y[118]; // @[G128Multiplay.scala 37:16:@2631.4]
  assign _T_659 = Z_9 ^ V_9; // @[G128Multiplay.scala 40:24:@2634.6]
  assign Z_10 = _T_656 ? _T_659 : Z_9; // @[G128Multiplay.scala 38:7:@2633.4]
  assign _T_660 = V_9[0]; // @[G128Multiplay.scala 45:18:@2640.4]
  assign _T_662 = _T_660 == 1'h0; // @[G128Multiplay.scala 45:22:@2641.4]
  assign _T_664 = V_9 >> 1'h1; // @[G128Multiplay.scala 48:24:@2643.6]
  assign _T_668 = _T_664 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2649.6]
  assign V_10 = _T_662 ? _T_664 : _T_668; // @[G128Multiplay.scala 46:7:@2642.4]
  assign _T_670 = io_y[117]; // @[G128Multiplay.scala 37:16:@2653.4]
  assign _T_673 = Z_10 ^ V_10; // @[G128Multiplay.scala 40:24:@2656.6]
  assign Z_11 = _T_670 ? _T_673 : Z_10; // @[G128Multiplay.scala 38:7:@2655.4]
  assign _T_674 = V_10[0]; // @[G128Multiplay.scala 45:18:@2662.4]
  assign _T_676 = _T_674 == 1'h0; // @[G128Multiplay.scala 45:22:@2663.4]
  assign _T_678 = V_10 >> 1'h1; // @[G128Multiplay.scala 48:24:@2665.6]
  assign _T_682 = _T_678 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2671.6]
  assign V_11 = _T_676 ? _T_678 : _T_682; // @[G128Multiplay.scala 46:7:@2664.4]
  assign _T_684 = io_y[116]; // @[G128Multiplay.scala 37:16:@2675.4]
  assign _T_687 = Z_11 ^ V_11; // @[G128Multiplay.scala 40:24:@2678.6]
  assign Z_12 = _T_684 ? _T_687 : Z_11; // @[G128Multiplay.scala 38:7:@2677.4]
  assign _T_688 = V_11[0]; // @[G128Multiplay.scala 45:18:@2684.4]
  assign _T_690 = _T_688 == 1'h0; // @[G128Multiplay.scala 45:22:@2685.4]
  assign _T_692 = V_11 >> 1'h1; // @[G128Multiplay.scala 48:24:@2687.6]
  assign _T_696 = _T_692 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2693.6]
  assign V_12 = _T_690 ? _T_692 : _T_696; // @[G128Multiplay.scala 46:7:@2686.4]
  assign _T_698 = io_y[115]; // @[G128Multiplay.scala 37:16:@2697.4]
  assign _T_701 = Z_12 ^ V_12; // @[G128Multiplay.scala 40:24:@2700.6]
  assign Z_13 = _T_698 ? _T_701 : Z_12; // @[G128Multiplay.scala 38:7:@2699.4]
  assign _T_702 = V_12[0]; // @[G128Multiplay.scala 45:18:@2706.4]
  assign _T_704 = _T_702 == 1'h0; // @[G128Multiplay.scala 45:22:@2707.4]
  assign _T_706 = V_12 >> 1'h1; // @[G128Multiplay.scala 48:24:@2709.6]
  assign _T_710 = _T_706 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2715.6]
  assign V_13 = _T_704 ? _T_706 : _T_710; // @[G128Multiplay.scala 46:7:@2708.4]
  assign _T_712 = io_y[114]; // @[G128Multiplay.scala 37:16:@2719.4]
  assign _T_715 = Z_13 ^ V_13; // @[G128Multiplay.scala 40:24:@2722.6]
  assign Z_14 = _T_712 ? _T_715 : Z_13; // @[G128Multiplay.scala 38:7:@2721.4]
  assign _T_716 = V_13[0]; // @[G128Multiplay.scala 45:18:@2728.4]
  assign _T_718 = _T_716 == 1'h0; // @[G128Multiplay.scala 45:22:@2729.4]
  assign _T_720 = V_13 >> 1'h1; // @[G128Multiplay.scala 48:24:@2731.6]
  assign _T_724 = _T_720 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2737.6]
  assign V_14 = _T_718 ? _T_720 : _T_724; // @[G128Multiplay.scala 46:7:@2730.4]
  assign _T_726 = io_y[113]; // @[G128Multiplay.scala 37:16:@2741.4]
  assign _T_729 = Z_14 ^ V_14; // @[G128Multiplay.scala 40:24:@2744.6]
  assign Z_15 = _T_726 ? _T_729 : Z_14; // @[G128Multiplay.scala 38:7:@2743.4]
  assign _T_730 = V_14[0]; // @[G128Multiplay.scala 45:18:@2750.4]
  assign _T_732 = _T_730 == 1'h0; // @[G128Multiplay.scala 45:22:@2751.4]
  assign _T_734 = V_14 >> 1'h1; // @[G128Multiplay.scala 48:24:@2753.6]
  assign _T_738 = _T_734 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2759.6]
  assign V_15 = _T_732 ? _T_734 : _T_738; // @[G128Multiplay.scala 46:7:@2752.4]
  assign _T_740 = io_y[112]; // @[G128Multiplay.scala 37:16:@2763.4]
  assign _T_743 = Z_15 ^ V_15; // @[G128Multiplay.scala 40:24:@2766.6]
  assign Z_16 = _T_740 ? _T_743 : Z_15; // @[G128Multiplay.scala 38:7:@2765.4]
  assign _T_744 = V_15[0]; // @[G128Multiplay.scala 45:18:@2772.4]
  assign _T_746 = _T_744 == 1'h0; // @[G128Multiplay.scala 45:22:@2773.4]
  assign _T_748 = V_15 >> 1'h1; // @[G128Multiplay.scala 48:24:@2775.6]
  assign _T_752 = _T_748 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2781.6]
  assign V_16 = _T_746 ? _T_748 : _T_752; // @[G128Multiplay.scala 46:7:@2774.4]
  assign _T_754 = io_y[111]; // @[G128Multiplay.scala 37:16:@2785.4]
  assign _T_757 = Z_16 ^ V_16; // @[G128Multiplay.scala 40:24:@2788.6]
  assign Z_17 = _T_754 ? _T_757 : Z_16; // @[G128Multiplay.scala 38:7:@2787.4]
  assign _T_758 = V_16[0]; // @[G128Multiplay.scala 45:18:@2794.4]
  assign _T_760 = _T_758 == 1'h0; // @[G128Multiplay.scala 45:22:@2795.4]
  assign _T_762 = V_16 >> 1'h1; // @[G128Multiplay.scala 48:24:@2797.6]
  assign _T_766 = _T_762 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2803.6]
  assign V_17 = _T_760 ? _T_762 : _T_766; // @[G128Multiplay.scala 46:7:@2796.4]
  assign _T_768 = io_y[110]; // @[G128Multiplay.scala 37:16:@2807.4]
  assign _T_771 = Z_17 ^ V_17; // @[G128Multiplay.scala 40:24:@2810.6]
  assign Z_18 = _T_768 ? _T_771 : Z_17; // @[G128Multiplay.scala 38:7:@2809.4]
  assign _T_772 = V_17[0]; // @[G128Multiplay.scala 45:18:@2816.4]
  assign _T_774 = _T_772 == 1'h0; // @[G128Multiplay.scala 45:22:@2817.4]
  assign _T_776 = V_17 >> 1'h1; // @[G128Multiplay.scala 48:24:@2819.6]
  assign _T_780 = _T_776 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2825.6]
  assign V_18 = _T_774 ? _T_776 : _T_780; // @[G128Multiplay.scala 46:7:@2818.4]
  assign _T_782 = io_y[109]; // @[G128Multiplay.scala 37:16:@2829.4]
  assign _T_785 = Z_18 ^ V_18; // @[G128Multiplay.scala 40:24:@2832.6]
  assign Z_19 = _T_782 ? _T_785 : Z_18; // @[G128Multiplay.scala 38:7:@2831.4]
  assign _T_786 = V_18[0]; // @[G128Multiplay.scala 45:18:@2838.4]
  assign _T_788 = _T_786 == 1'h0; // @[G128Multiplay.scala 45:22:@2839.4]
  assign _T_790 = V_18 >> 1'h1; // @[G128Multiplay.scala 48:24:@2841.6]
  assign _T_794 = _T_790 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2847.6]
  assign V_19 = _T_788 ? _T_790 : _T_794; // @[G128Multiplay.scala 46:7:@2840.4]
  assign _T_796 = io_y[108]; // @[G128Multiplay.scala 37:16:@2851.4]
  assign _T_799 = Z_19 ^ V_19; // @[G128Multiplay.scala 40:24:@2854.6]
  assign Z_20 = _T_796 ? _T_799 : Z_19; // @[G128Multiplay.scala 38:7:@2853.4]
  assign _T_800 = V_19[0]; // @[G128Multiplay.scala 45:18:@2860.4]
  assign _T_802 = _T_800 == 1'h0; // @[G128Multiplay.scala 45:22:@2861.4]
  assign _T_804 = V_19 >> 1'h1; // @[G128Multiplay.scala 48:24:@2863.6]
  assign _T_808 = _T_804 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2869.6]
  assign V_20 = _T_802 ? _T_804 : _T_808; // @[G128Multiplay.scala 46:7:@2862.4]
  assign _T_810 = io_y[107]; // @[G128Multiplay.scala 37:16:@2873.4]
  assign _T_813 = Z_20 ^ V_20; // @[G128Multiplay.scala 40:24:@2876.6]
  assign Z_21 = _T_810 ? _T_813 : Z_20; // @[G128Multiplay.scala 38:7:@2875.4]
  assign _T_814 = V_20[0]; // @[G128Multiplay.scala 45:18:@2882.4]
  assign _T_816 = _T_814 == 1'h0; // @[G128Multiplay.scala 45:22:@2883.4]
  assign _T_818 = V_20 >> 1'h1; // @[G128Multiplay.scala 48:24:@2885.6]
  assign _T_822 = _T_818 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2891.6]
  assign V_21 = _T_816 ? _T_818 : _T_822; // @[G128Multiplay.scala 46:7:@2884.4]
  assign _T_824 = io_y[106]; // @[G128Multiplay.scala 37:16:@2895.4]
  assign _T_827 = Z_21 ^ V_21; // @[G128Multiplay.scala 40:24:@2898.6]
  assign Z_22 = _T_824 ? _T_827 : Z_21; // @[G128Multiplay.scala 38:7:@2897.4]
  assign _T_828 = V_21[0]; // @[G128Multiplay.scala 45:18:@2904.4]
  assign _T_830 = _T_828 == 1'h0; // @[G128Multiplay.scala 45:22:@2905.4]
  assign _T_832 = V_21 >> 1'h1; // @[G128Multiplay.scala 48:24:@2907.6]
  assign _T_836 = _T_832 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2913.6]
  assign V_22 = _T_830 ? _T_832 : _T_836; // @[G128Multiplay.scala 46:7:@2906.4]
  assign _T_838 = io_y[105]; // @[G128Multiplay.scala 37:16:@2917.4]
  assign _T_841 = Z_22 ^ V_22; // @[G128Multiplay.scala 40:24:@2920.6]
  assign Z_23 = _T_838 ? _T_841 : Z_22; // @[G128Multiplay.scala 38:7:@2919.4]
  assign _T_842 = V_22[0]; // @[G128Multiplay.scala 45:18:@2926.4]
  assign _T_844 = _T_842 == 1'h0; // @[G128Multiplay.scala 45:22:@2927.4]
  assign _T_846 = V_22 >> 1'h1; // @[G128Multiplay.scala 48:24:@2929.6]
  assign _T_850 = _T_846 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2935.6]
  assign V_23 = _T_844 ? _T_846 : _T_850; // @[G128Multiplay.scala 46:7:@2928.4]
  assign _T_852 = io_y[104]; // @[G128Multiplay.scala 37:16:@2939.4]
  assign _T_855 = Z_23 ^ V_23; // @[G128Multiplay.scala 40:24:@2942.6]
  assign Z_24 = _T_852 ? _T_855 : Z_23; // @[G128Multiplay.scala 38:7:@2941.4]
  assign _T_856 = V_23[0]; // @[G128Multiplay.scala 45:18:@2948.4]
  assign _T_858 = _T_856 == 1'h0; // @[G128Multiplay.scala 45:22:@2949.4]
  assign _T_860 = V_23 >> 1'h1; // @[G128Multiplay.scala 48:24:@2951.6]
  assign _T_864 = _T_860 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2957.6]
  assign V_24 = _T_858 ? _T_860 : _T_864; // @[G128Multiplay.scala 46:7:@2950.4]
  assign _T_866 = io_y[103]; // @[G128Multiplay.scala 37:16:@2961.4]
  assign _T_869 = Z_24 ^ V_24; // @[G128Multiplay.scala 40:24:@2964.6]
  assign Z_25 = _T_866 ? _T_869 : Z_24; // @[G128Multiplay.scala 38:7:@2963.4]
  assign _T_870 = V_24[0]; // @[G128Multiplay.scala 45:18:@2970.4]
  assign _T_872 = _T_870 == 1'h0; // @[G128Multiplay.scala 45:22:@2971.4]
  assign _T_874 = V_24 >> 1'h1; // @[G128Multiplay.scala 48:24:@2973.6]
  assign _T_878 = _T_874 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@2979.6]
  assign V_25 = _T_872 ? _T_874 : _T_878; // @[G128Multiplay.scala 46:7:@2972.4]
  assign _T_880 = io_y[102]; // @[G128Multiplay.scala 37:16:@2983.4]
  assign _T_883 = Z_25 ^ V_25; // @[G128Multiplay.scala 40:24:@2986.6]
  assign Z_26 = _T_880 ? _T_883 : Z_25; // @[G128Multiplay.scala 38:7:@2985.4]
  assign _T_884 = V_25[0]; // @[G128Multiplay.scala 45:18:@2992.4]
  assign _T_886 = _T_884 == 1'h0; // @[G128Multiplay.scala 45:22:@2993.4]
  assign _T_888 = V_25 >> 1'h1; // @[G128Multiplay.scala 48:24:@2995.6]
  assign _T_892 = _T_888 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3001.6]
  assign V_26 = _T_886 ? _T_888 : _T_892; // @[G128Multiplay.scala 46:7:@2994.4]
  assign _T_894 = io_y[101]; // @[G128Multiplay.scala 37:16:@3005.4]
  assign _T_897 = Z_26 ^ V_26; // @[G128Multiplay.scala 40:24:@3008.6]
  assign Z_27 = _T_894 ? _T_897 : Z_26; // @[G128Multiplay.scala 38:7:@3007.4]
  assign _T_898 = V_26[0]; // @[G128Multiplay.scala 45:18:@3014.4]
  assign _T_900 = _T_898 == 1'h0; // @[G128Multiplay.scala 45:22:@3015.4]
  assign _T_902 = V_26 >> 1'h1; // @[G128Multiplay.scala 48:24:@3017.6]
  assign _T_906 = _T_902 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3023.6]
  assign V_27 = _T_900 ? _T_902 : _T_906; // @[G128Multiplay.scala 46:7:@3016.4]
  assign _T_908 = io_y[100]; // @[G128Multiplay.scala 37:16:@3027.4]
  assign _T_911 = Z_27 ^ V_27; // @[G128Multiplay.scala 40:24:@3030.6]
  assign Z_28 = _T_908 ? _T_911 : Z_27; // @[G128Multiplay.scala 38:7:@3029.4]
  assign _T_912 = V_27[0]; // @[G128Multiplay.scala 45:18:@3036.4]
  assign _T_914 = _T_912 == 1'h0; // @[G128Multiplay.scala 45:22:@3037.4]
  assign _T_916 = V_27 >> 1'h1; // @[G128Multiplay.scala 48:24:@3039.6]
  assign _T_920 = _T_916 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3045.6]
  assign V_28 = _T_914 ? _T_916 : _T_920; // @[G128Multiplay.scala 46:7:@3038.4]
  assign _T_922 = io_y[99]; // @[G128Multiplay.scala 37:16:@3049.4]
  assign _T_925 = Z_28 ^ V_28; // @[G128Multiplay.scala 40:24:@3052.6]
  assign Z_29 = _T_922 ? _T_925 : Z_28; // @[G128Multiplay.scala 38:7:@3051.4]
  assign _T_926 = V_28[0]; // @[G128Multiplay.scala 45:18:@3058.4]
  assign _T_928 = _T_926 == 1'h0; // @[G128Multiplay.scala 45:22:@3059.4]
  assign _T_930 = V_28 >> 1'h1; // @[G128Multiplay.scala 48:24:@3061.6]
  assign _T_934 = _T_930 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3067.6]
  assign V_29 = _T_928 ? _T_930 : _T_934; // @[G128Multiplay.scala 46:7:@3060.4]
  assign _T_936 = io_y[98]; // @[G128Multiplay.scala 37:16:@3071.4]
  assign _T_939 = Z_29 ^ V_29; // @[G128Multiplay.scala 40:24:@3074.6]
  assign Z_30 = _T_936 ? _T_939 : Z_29; // @[G128Multiplay.scala 38:7:@3073.4]
  assign _T_940 = V_29[0]; // @[G128Multiplay.scala 45:18:@3080.4]
  assign _T_942 = _T_940 == 1'h0; // @[G128Multiplay.scala 45:22:@3081.4]
  assign _T_944 = V_29 >> 1'h1; // @[G128Multiplay.scala 48:24:@3083.6]
  assign _T_948 = _T_944 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3089.6]
  assign V_30 = _T_942 ? _T_944 : _T_948; // @[G128Multiplay.scala 46:7:@3082.4]
  assign _T_950 = io_y[97]; // @[G128Multiplay.scala 37:16:@3093.4]
  assign _T_953 = Z_30 ^ V_30; // @[G128Multiplay.scala 40:24:@3096.6]
  assign Z_31 = _T_950 ? _T_953 : Z_30; // @[G128Multiplay.scala 38:7:@3095.4]
  assign _T_954 = V_30[0]; // @[G128Multiplay.scala 45:18:@3102.4]
  assign _T_956 = _T_954 == 1'h0; // @[G128Multiplay.scala 45:22:@3103.4]
  assign _T_958 = V_30 >> 1'h1; // @[G128Multiplay.scala 48:24:@3105.6]
  assign _T_962 = _T_958 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3111.6]
  assign V_31 = _T_956 ? _T_958 : _T_962; // @[G128Multiplay.scala 46:7:@3104.4]
  assign _T_964 = io_y[96]; // @[G128Multiplay.scala 37:16:@3115.4]
  assign _T_967 = Z_31 ^ V_31; // @[G128Multiplay.scala 40:24:@3118.6]
  assign Z_32 = _T_964 ? _T_967 : Z_31; // @[G128Multiplay.scala 38:7:@3117.4]
  assign _T_968 = V_31[0]; // @[G128Multiplay.scala 45:18:@3124.4]
  assign _T_970 = _T_968 == 1'h0; // @[G128Multiplay.scala 45:22:@3125.4]
  assign _T_972 = V_31 >> 1'h1; // @[G128Multiplay.scala 48:24:@3127.6]
  assign _T_976 = _T_972 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3133.6]
  assign V_32 = _T_970 ? _T_972 : _T_976; // @[G128Multiplay.scala 46:7:@3126.4]
  assign _T_978 = io_y[95]; // @[G128Multiplay.scala 37:16:@3137.4]
  assign _T_981 = Z_32 ^ V_32; // @[G128Multiplay.scala 40:24:@3140.6]
  assign Z_33 = _T_978 ? _T_981 : Z_32; // @[G128Multiplay.scala 38:7:@3139.4]
  assign _T_982 = V_32[0]; // @[G128Multiplay.scala 45:18:@3146.4]
  assign _T_984 = _T_982 == 1'h0; // @[G128Multiplay.scala 45:22:@3147.4]
  assign _T_986 = V_32 >> 1'h1; // @[G128Multiplay.scala 48:24:@3149.6]
  assign _T_990 = _T_986 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3155.6]
  assign V_33 = _T_984 ? _T_986 : _T_990; // @[G128Multiplay.scala 46:7:@3148.4]
  assign _T_992 = io_y[94]; // @[G128Multiplay.scala 37:16:@3159.4]
  assign _T_995 = Z_33 ^ V_33; // @[G128Multiplay.scala 40:24:@3162.6]
  assign Z_34 = _T_992 ? _T_995 : Z_33; // @[G128Multiplay.scala 38:7:@3161.4]
  assign _T_996 = V_33[0]; // @[G128Multiplay.scala 45:18:@3168.4]
  assign _T_998 = _T_996 == 1'h0; // @[G128Multiplay.scala 45:22:@3169.4]
  assign _T_1000 = V_33 >> 1'h1; // @[G128Multiplay.scala 48:24:@3171.6]
  assign _T_1004 = _T_1000 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3177.6]
  assign V_34 = _T_998 ? _T_1000 : _T_1004; // @[G128Multiplay.scala 46:7:@3170.4]
  assign _T_1006 = io_y[93]; // @[G128Multiplay.scala 37:16:@3181.4]
  assign _T_1009 = Z_34 ^ V_34; // @[G128Multiplay.scala 40:24:@3184.6]
  assign Z_35 = _T_1006 ? _T_1009 : Z_34; // @[G128Multiplay.scala 38:7:@3183.4]
  assign _T_1010 = V_34[0]; // @[G128Multiplay.scala 45:18:@3190.4]
  assign _T_1012 = _T_1010 == 1'h0; // @[G128Multiplay.scala 45:22:@3191.4]
  assign _T_1014 = V_34 >> 1'h1; // @[G128Multiplay.scala 48:24:@3193.6]
  assign _T_1018 = _T_1014 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3199.6]
  assign V_35 = _T_1012 ? _T_1014 : _T_1018; // @[G128Multiplay.scala 46:7:@3192.4]
  assign _T_1020 = io_y[92]; // @[G128Multiplay.scala 37:16:@3203.4]
  assign _T_1023 = Z_35 ^ V_35; // @[G128Multiplay.scala 40:24:@3206.6]
  assign Z_36 = _T_1020 ? _T_1023 : Z_35; // @[G128Multiplay.scala 38:7:@3205.4]
  assign _T_1024 = V_35[0]; // @[G128Multiplay.scala 45:18:@3212.4]
  assign _T_1026 = _T_1024 == 1'h0; // @[G128Multiplay.scala 45:22:@3213.4]
  assign _T_1028 = V_35 >> 1'h1; // @[G128Multiplay.scala 48:24:@3215.6]
  assign _T_1032 = _T_1028 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3221.6]
  assign V_36 = _T_1026 ? _T_1028 : _T_1032; // @[G128Multiplay.scala 46:7:@3214.4]
  assign _T_1034 = io_y[91]; // @[G128Multiplay.scala 37:16:@3225.4]
  assign _T_1037 = Z_36 ^ V_36; // @[G128Multiplay.scala 40:24:@3228.6]
  assign Z_37 = _T_1034 ? _T_1037 : Z_36; // @[G128Multiplay.scala 38:7:@3227.4]
  assign _T_1038 = V_36[0]; // @[G128Multiplay.scala 45:18:@3234.4]
  assign _T_1040 = _T_1038 == 1'h0; // @[G128Multiplay.scala 45:22:@3235.4]
  assign _T_1042 = V_36 >> 1'h1; // @[G128Multiplay.scala 48:24:@3237.6]
  assign _T_1046 = _T_1042 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3243.6]
  assign V_37 = _T_1040 ? _T_1042 : _T_1046; // @[G128Multiplay.scala 46:7:@3236.4]
  assign _T_1048 = io_y[90]; // @[G128Multiplay.scala 37:16:@3247.4]
  assign _T_1051 = Z_37 ^ V_37; // @[G128Multiplay.scala 40:24:@3250.6]
  assign Z_38 = _T_1048 ? _T_1051 : Z_37; // @[G128Multiplay.scala 38:7:@3249.4]
  assign _T_1052 = V_37[0]; // @[G128Multiplay.scala 45:18:@3256.4]
  assign _T_1054 = _T_1052 == 1'h0; // @[G128Multiplay.scala 45:22:@3257.4]
  assign _T_1056 = V_37 >> 1'h1; // @[G128Multiplay.scala 48:24:@3259.6]
  assign _T_1060 = _T_1056 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3265.6]
  assign V_38 = _T_1054 ? _T_1056 : _T_1060; // @[G128Multiplay.scala 46:7:@3258.4]
  assign _T_1062 = io_y[89]; // @[G128Multiplay.scala 37:16:@3269.4]
  assign _T_1065 = Z_38 ^ V_38; // @[G128Multiplay.scala 40:24:@3272.6]
  assign Z_39 = _T_1062 ? _T_1065 : Z_38; // @[G128Multiplay.scala 38:7:@3271.4]
  assign _T_1066 = V_38[0]; // @[G128Multiplay.scala 45:18:@3278.4]
  assign _T_1068 = _T_1066 == 1'h0; // @[G128Multiplay.scala 45:22:@3279.4]
  assign _T_1070 = V_38 >> 1'h1; // @[G128Multiplay.scala 48:24:@3281.6]
  assign _T_1074 = _T_1070 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3287.6]
  assign V_39 = _T_1068 ? _T_1070 : _T_1074; // @[G128Multiplay.scala 46:7:@3280.4]
  assign _T_1076 = io_y[88]; // @[G128Multiplay.scala 37:16:@3291.4]
  assign _T_1079 = Z_39 ^ V_39; // @[G128Multiplay.scala 40:24:@3294.6]
  assign Z_40 = _T_1076 ? _T_1079 : Z_39; // @[G128Multiplay.scala 38:7:@3293.4]
  assign _T_1080 = V_39[0]; // @[G128Multiplay.scala 45:18:@3300.4]
  assign _T_1082 = _T_1080 == 1'h0; // @[G128Multiplay.scala 45:22:@3301.4]
  assign _T_1084 = V_39 >> 1'h1; // @[G128Multiplay.scala 48:24:@3303.6]
  assign _T_1088 = _T_1084 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3309.6]
  assign V_40 = _T_1082 ? _T_1084 : _T_1088; // @[G128Multiplay.scala 46:7:@3302.4]
  assign _T_1090 = io_y[87]; // @[G128Multiplay.scala 37:16:@3313.4]
  assign _T_1093 = Z_40 ^ V_40; // @[G128Multiplay.scala 40:24:@3316.6]
  assign Z_41 = _T_1090 ? _T_1093 : Z_40; // @[G128Multiplay.scala 38:7:@3315.4]
  assign _T_1094 = V_40[0]; // @[G128Multiplay.scala 45:18:@3322.4]
  assign _T_1096 = _T_1094 == 1'h0; // @[G128Multiplay.scala 45:22:@3323.4]
  assign _T_1098 = V_40 >> 1'h1; // @[G128Multiplay.scala 48:24:@3325.6]
  assign _T_1102 = _T_1098 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3331.6]
  assign V_41 = _T_1096 ? _T_1098 : _T_1102; // @[G128Multiplay.scala 46:7:@3324.4]
  assign _T_1104 = io_y[86]; // @[G128Multiplay.scala 37:16:@3335.4]
  assign _T_1107 = Z_41 ^ V_41; // @[G128Multiplay.scala 40:24:@3338.6]
  assign Z_42 = _T_1104 ? _T_1107 : Z_41; // @[G128Multiplay.scala 38:7:@3337.4]
  assign _T_1108 = V_41[0]; // @[G128Multiplay.scala 45:18:@3344.4]
  assign _T_1110 = _T_1108 == 1'h0; // @[G128Multiplay.scala 45:22:@3345.4]
  assign _T_1112 = V_41 >> 1'h1; // @[G128Multiplay.scala 48:24:@3347.6]
  assign _T_1116 = _T_1112 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3353.6]
  assign V_42 = _T_1110 ? _T_1112 : _T_1116; // @[G128Multiplay.scala 46:7:@3346.4]
  assign _T_1118 = io_y[85]; // @[G128Multiplay.scala 37:16:@3357.4]
  assign _T_1121 = Z_42 ^ V_42; // @[G128Multiplay.scala 40:24:@3360.6]
  assign Z_43 = _T_1118 ? _T_1121 : Z_42; // @[G128Multiplay.scala 38:7:@3359.4]
  assign _T_1122 = V_42[0]; // @[G128Multiplay.scala 45:18:@3366.4]
  assign _T_1124 = _T_1122 == 1'h0; // @[G128Multiplay.scala 45:22:@3367.4]
  assign _T_1126 = V_42 >> 1'h1; // @[G128Multiplay.scala 48:24:@3369.6]
  assign _T_1130 = _T_1126 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3375.6]
  assign V_43 = _T_1124 ? _T_1126 : _T_1130; // @[G128Multiplay.scala 46:7:@3368.4]
  assign _T_1132 = io_y[84]; // @[G128Multiplay.scala 37:16:@3379.4]
  assign _T_1135 = Z_43 ^ V_43; // @[G128Multiplay.scala 40:24:@3382.6]
  assign Z_44 = _T_1132 ? _T_1135 : Z_43; // @[G128Multiplay.scala 38:7:@3381.4]
  assign _T_1136 = V_43[0]; // @[G128Multiplay.scala 45:18:@3388.4]
  assign _T_1138 = _T_1136 == 1'h0; // @[G128Multiplay.scala 45:22:@3389.4]
  assign _T_1140 = V_43 >> 1'h1; // @[G128Multiplay.scala 48:24:@3391.6]
  assign _T_1144 = _T_1140 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3397.6]
  assign V_44 = _T_1138 ? _T_1140 : _T_1144; // @[G128Multiplay.scala 46:7:@3390.4]
  assign _T_1146 = io_y[83]; // @[G128Multiplay.scala 37:16:@3401.4]
  assign _T_1149 = Z_44 ^ V_44; // @[G128Multiplay.scala 40:24:@3404.6]
  assign Z_45 = _T_1146 ? _T_1149 : Z_44; // @[G128Multiplay.scala 38:7:@3403.4]
  assign _T_1150 = V_44[0]; // @[G128Multiplay.scala 45:18:@3410.4]
  assign _T_1152 = _T_1150 == 1'h0; // @[G128Multiplay.scala 45:22:@3411.4]
  assign _T_1154 = V_44 >> 1'h1; // @[G128Multiplay.scala 48:24:@3413.6]
  assign _T_1158 = _T_1154 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3419.6]
  assign V_45 = _T_1152 ? _T_1154 : _T_1158; // @[G128Multiplay.scala 46:7:@3412.4]
  assign _T_1160 = io_y[82]; // @[G128Multiplay.scala 37:16:@3423.4]
  assign _T_1163 = Z_45 ^ V_45; // @[G128Multiplay.scala 40:24:@3426.6]
  assign Z_46 = _T_1160 ? _T_1163 : Z_45; // @[G128Multiplay.scala 38:7:@3425.4]
  assign _T_1164 = V_45[0]; // @[G128Multiplay.scala 45:18:@3432.4]
  assign _T_1166 = _T_1164 == 1'h0; // @[G128Multiplay.scala 45:22:@3433.4]
  assign _T_1168 = V_45 >> 1'h1; // @[G128Multiplay.scala 48:24:@3435.6]
  assign _T_1172 = _T_1168 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3441.6]
  assign V_46 = _T_1166 ? _T_1168 : _T_1172; // @[G128Multiplay.scala 46:7:@3434.4]
  assign _T_1174 = io_y[81]; // @[G128Multiplay.scala 37:16:@3445.4]
  assign _T_1177 = Z_46 ^ V_46; // @[G128Multiplay.scala 40:24:@3448.6]
  assign Z_47 = _T_1174 ? _T_1177 : Z_46; // @[G128Multiplay.scala 38:7:@3447.4]
  assign _T_1178 = V_46[0]; // @[G128Multiplay.scala 45:18:@3454.4]
  assign _T_1180 = _T_1178 == 1'h0; // @[G128Multiplay.scala 45:22:@3455.4]
  assign _T_1182 = V_46 >> 1'h1; // @[G128Multiplay.scala 48:24:@3457.6]
  assign _T_1186 = _T_1182 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3463.6]
  assign V_47 = _T_1180 ? _T_1182 : _T_1186; // @[G128Multiplay.scala 46:7:@3456.4]
  assign _T_1188 = io_y[80]; // @[G128Multiplay.scala 37:16:@3467.4]
  assign _T_1191 = Z_47 ^ V_47; // @[G128Multiplay.scala 40:24:@3470.6]
  assign Z_48 = _T_1188 ? _T_1191 : Z_47; // @[G128Multiplay.scala 38:7:@3469.4]
  assign _T_1192 = V_47[0]; // @[G128Multiplay.scala 45:18:@3476.4]
  assign _T_1194 = _T_1192 == 1'h0; // @[G128Multiplay.scala 45:22:@3477.4]
  assign _T_1196 = V_47 >> 1'h1; // @[G128Multiplay.scala 48:24:@3479.6]
  assign _T_1200 = _T_1196 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3485.6]
  assign V_48 = _T_1194 ? _T_1196 : _T_1200; // @[G128Multiplay.scala 46:7:@3478.4]
  assign _T_1202 = io_y[79]; // @[G128Multiplay.scala 37:16:@3489.4]
  assign _T_1205 = Z_48 ^ V_48; // @[G128Multiplay.scala 40:24:@3492.6]
  assign Z_49 = _T_1202 ? _T_1205 : Z_48; // @[G128Multiplay.scala 38:7:@3491.4]
  assign _T_1206 = V_48[0]; // @[G128Multiplay.scala 45:18:@3498.4]
  assign _T_1208 = _T_1206 == 1'h0; // @[G128Multiplay.scala 45:22:@3499.4]
  assign _T_1210 = V_48 >> 1'h1; // @[G128Multiplay.scala 48:24:@3501.6]
  assign _T_1214 = _T_1210 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3507.6]
  assign V_49 = _T_1208 ? _T_1210 : _T_1214; // @[G128Multiplay.scala 46:7:@3500.4]
  assign _T_1216 = io_y[78]; // @[G128Multiplay.scala 37:16:@3511.4]
  assign _T_1219 = Z_49 ^ V_49; // @[G128Multiplay.scala 40:24:@3514.6]
  assign Z_50 = _T_1216 ? _T_1219 : Z_49; // @[G128Multiplay.scala 38:7:@3513.4]
  assign _T_1220 = V_49[0]; // @[G128Multiplay.scala 45:18:@3520.4]
  assign _T_1222 = _T_1220 == 1'h0; // @[G128Multiplay.scala 45:22:@3521.4]
  assign _T_1224 = V_49 >> 1'h1; // @[G128Multiplay.scala 48:24:@3523.6]
  assign _T_1228 = _T_1224 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3529.6]
  assign V_50 = _T_1222 ? _T_1224 : _T_1228; // @[G128Multiplay.scala 46:7:@3522.4]
  assign _T_1230 = io_y[77]; // @[G128Multiplay.scala 37:16:@3533.4]
  assign _T_1233 = Z_50 ^ V_50; // @[G128Multiplay.scala 40:24:@3536.6]
  assign Z_51 = _T_1230 ? _T_1233 : Z_50; // @[G128Multiplay.scala 38:7:@3535.4]
  assign _T_1234 = V_50[0]; // @[G128Multiplay.scala 45:18:@3542.4]
  assign _T_1236 = _T_1234 == 1'h0; // @[G128Multiplay.scala 45:22:@3543.4]
  assign _T_1238 = V_50 >> 1'h1; // @[G128Multiplay.scala 48:24:@3545.6]
  assign _T_1242 = _T_1238 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3551.6]
  assign V_51 = _T_1236 ? _T_1238 : _T_1242; // @[G128Multiplay.scala 46:7:@3544.4]
  assign _T_1244 = io_y[76]; // @[G128Multiplay.scala 37:16:@3555.4]
  assign _T_1247 = Z_51 ^ V_51; // @[G128Multiplay.scala 40:24:@3558.6]
  assign Z_52 = _T_1244 ? _T_1247 : Z_51; // @[G128Multiplay.scala 38:7:@3557.4]
  assign _T_1248 = V_51[0]; // @[G128Multiplay.scala 45:18:@3564.4]
  assign _T_1250 = _T_1248 == 1'h0; // @[G128Multiplay.scala 45:22:@3565.4]
  assign _T_1252 = V_51 >> 1'h1; // @[G128Multiplay.scala 48:24:@3567.6]
  assign _T_1256 = _T_1252 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3573.6]
  assign V_52 = _T_1250 ? _T_1252 : _T_1256; // @[G128Multiplay.scala 46:7:@3566.4]
  assign _T_1258 = io_y[75]; // @[G128Multiplay.scala 37:16:@3577.4]
  assign _T_1261 = Z_52 ^ V_52; // @[G128Multiplay.scala 40:24:@3580.6]
  assign Z_53 = _T_1258 ? _T_1261 : Z_52; // @[G128Multiplay.scala 38:7:@3579.4]
  assign _T_1262 = V_52[0]; // @[G128Multiplay.scala 45:18:@3586.4]
  assign _T_1264 = _T_1262 == 1'h0; // @[G128Multiplay.scala 45:22:@3587.4]
  assign _T_1266 = V_52 >> 1'h1; // @[G128Multiplay.scala 48:24:@3589.6]
  assign _T_1270 = _T_1266 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3595.6]
  assign V_53 = _T_1264 ? _T_1266 : _T_1270; // @[G128Multiplay.scala 46:7:@3588.4]
  assign _T_1272 = io_y[74]; // @[G128Multiplay.scala 37:16:@3599.4]
  assign _T_1275 = Z_53 ^ V_53; // @[G128Multiplay.scala 40:24:@3602.6]
  assign Z_54 = _T_1272 ? _T_1275 : Z_53; // @[G128Multiplay.scala 38:7:@3601.4]
  assign _T_1276 = V_53[0]; // @[G128Multiplay.scala 45:18:@3608.4]
  assign _T_1278 = _T_1276 == 1'h0; // @[G128Multiplay.scala 45:22:@3609.4]
  assign _T_1280 = V_53 >> 1'h1; // @[G128Multiplay.scala 48:24:@3611.6]
  assign _T_1284 = _T_1280 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3617.6]
  assign V_54 = _T_1278 ? _T_1280 : _T_1284; // @[G128Multiplay.scala 46:7:@3610.4]
  assign _T_1286 = io_y[73]; // @[G128Multiplay.scala 37:16:@3621.4]
  assign _T_1289 = Z_54 ^ V_54; // @[G128Multiplay.scala 40:24:@3624.6]
  assign Z_55 = _T_1286 ? _T_1289 : Z_54; // @[G128Multiplay.scala 38:7:@3623.4]
  assign _T_1290 = V_54[0]; // @[G128Multiplay.scala 45:18:@3630.4]
  assign _T_1292 = _T_1290 == 1'h0; // @[G128Multiplay.scala 45:22:@3631.4]
  assign _T_1294 = V_54 >> 1'h1; // @[G128Multiplay.scala 48:24:@3633.6]
  assign _T_1298 = _T_1294 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3639.6]
  assign V_55 = _T_1292 ? _T_1294 : _T_1298; // @[G128Multiplay.scala 46:7:@3632.4]
  assign _T_1300 = io_y[72]; // @[G128Multiplay.scala 37:16:@3643.4]
  assign _T_1303 = Z_55 ^ V_55; // @[G128Multiplay.scala 40:24:@3646.6]
  assign Z_56 = _T_1300 ? _T_1303 : Z_55; // @[G128Multiplay.scala 38:7:@3645.4]
  assign _T_1304 = V_55[0]; // @[G128Multiplay.scala 45:18:@3652.4]
  assign _T_1306 = _T_1304 == 1'h0; // @[G128Multiplay.scala 45:22:@3653.4]
  assign _T_1308 = V_55 >> 1'h1; // @[G128Multiplay.scala 48:24:@3655.6]
  assign _T_1312 = _T_1308 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3661.6]
  assign V_56 = _T_1306 ? _T_1308 : _T_1312; // @[G128Multiplay.scala 46:7:@3654.4]
  assign _T_1314 = io_y[71]; // @[G128Multiplay.scala 37:16:@3665.4]
  assign _T_1317 = Z_56 ^ V_56; // @[G128Multiplay.scala 40:24:@3668.6]
  assign Z_57 = _T_1314 ? _T_1317 : Z_56; // @[G128Multiplay.scala 38:7:@3667.4]
  assign _T_1318 = V_56[0]; // @[G128Multiplay.scala 45:18:@3674.4]
  assign _T_1320 = _T_1318 == 1'h0; // @[G128Multiplay.scala 45:22:@3675.4]
  assign _T_1322 = V_56 >> 1'h1; // @[G128Multiplay.scala 48:24:@3677.6]
  assign _T_1326 = _T_1322 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3683.6]
  assign V_57 = _T_1320 ? _T_1322 : _T_1326; // @[G128Multiplay.scala 46:7:@3676.4]
  assign _T_1328 = io_y[70]; // @[G128Multiplay.scala 37:16:@3687.4]
  assign _T_1331 = Z_57 ^ V_57; // @[G128Multiplay.scala 40:24:@3690.6]
  assign Z_58 = _T_1328 ? _T_1331 : Z_57; // @[G128Multiplay.scala 38:7:@3689.4]
  assign _T_1332 = V_57[0]; // @[G128Multiplay.scala 45:18:@3696.4]
  assign _T_1334 = _T_1332 == 1'h0; // @[G128Multiplay.scala 45:22:@3697.4]
  assign _T_1336 = V_57 >> 1'h1; // @[G128Multiplay.scala 48:24:@3699.6]
  assign _T_1340 = _T_1336 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3705.6]
  assign V_58 = _T_1334 ? _T_1336 : _T_1340; // @[G128Multiplay.scala 46:7:@3698.4]
  assign _T_1342 = io_y[69]; // @[G128Multiplay.scala 37:16:@3709.4]
  assign _T_1345 = Z_58 ^ V_58; // @[G128Multiplay.scala 40:24:@3712.6]
  assign Z_59 = _T_1342 ? _T_1345 : Z_58; // @[G128Multiplay.scala 38:7:@3711.4]
  assign _T_1346 = V_58[0]; // @[G128Multiplay.scala 45:18:@3718.4]
  assign _T_1348 = _T_1346 == 1'h0; // @[G128Multiplay.scala 45:22:@3719.4]
  assign _T_1350 = V_58 >> 1'h1; // @[G128Multiplay.scala 48:24:@3721.6]
  assign _T_1354 = _T_1350 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3727.6]
  assign V_59 = _T_1348 ? _T_1350 : _T_1354; // @[G128Multiplay.scala 46:7:@3720.4]
  assign _T_1356 = io_y[68]; // @[G128Multiplay.scala 37:16:@3731.4]
  assign _T_1359 = Z_59 ^ V_59; // @[G128Multiplay.scala 40:24:@3734.6]
  assign Z_60 = _T_1356 ? _T_1359 : Z_59; // @[G128Multiplay.scala 38:7:@3733.4]
  assign _T_1360 = V_59[0]; // @[G128Multiplay.scala 45:18:@3740.4]
  assign _T_1362 = _T_1360 == 1'h0; // @[G128Multiplay.scala 45:22:@3741.4]
  assign _T_1364 = V_59 >> 1'h1; // @[G128Multiplay.scala 48:24:@3743.6]
  assign _T_1368 = _T_1364 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3749.6]
  assign V_60 = _T_1362 ? _T_1364 : _T_1368; // @[G128Multiplay.scala 46:7:@3742.4]
  assign _T_1370 = io_y[67]; // @[G128Multiplay.scala 37:16:@3753.4]
  assign _T_1373 = Z_60 ^ V_60; // @[G128Multiplay.scala 40:24:@3756.6]
  assign Z_61 = _T_1370 ? _T_1373 : Z_60; // @[G128Multiplay.scala 38:7:@3755.4]
  assign _T_1374 = V_60[0]; // @[G128Multiplay.scala 45:18:@3762.4]
  assign _T_1376 = _T_1374 == 1'h0; // @[G128Multiplay.scala 45:22:@3763.4]
  assign _T_1378 = V_60 >> 1'h1; // @[G128Multiplay.scala 48:24:@3765.6]
  assign _T_1382 = _T_1378 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3771.6]
  assign V_61 = _T_1376 ? _T_1378 : _T_1382; // @[G128Multiplay.scala 46:7:@3764.4]
  assign _T_1384 = io_y[66]; // @[G128Multiplay.scala 37:16:@3775.4]
  assign _T_1387 = Z_61 ^ V_61; // @[G128Multiplay.scala 40:24:@3778.6]
  assign Z_62 = _T_1384 ? _T_1387 : Z_61; // @[G128Multiplay.scala 38:7:@3777.4]
  assign _T_1388 = V_61[0]; // @[G128Multiplay.scala 45:18:@3784.4]
  assign _T_1390 = _T_1388 == 1'h0; // @[G128Multiplay.scala 45:22:@3785.4]
  assign _T_1392 = V_61 >> 1'h1; // @[G128Multiplay.scala 48:24:@3787.6]
  assign _T_1396 = _T_1392 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3793.6]
  assign V_62 = _T_1390 ? _T_1392 : _T_1396; // @[G128Multiplay.scala 46:7:@3786.4]
  assign _T_1398 = io_y[65]; // @[G128Multiplay.scala 37:16:@3797.4]
  assign _T_1401 = Z_62 ^ V_62; // @[G128Multiplay.scala 40:24:@3800.6]
  assign Z_63 = _T_1398 ? _T_1401 : Z_62; // @[G128Multiplay.scala 38:7:@3799.4]
  assign _T_1402 = V_62[0]; // @[G128Multiplay.scala 45:18:@3806.4]
  assign _T_1404 = _T_1402 == 1'h0; // @[G128Multiplay.scala 45:22:@3807.4]
  assign _T_1406 = V_62 >> 1'h1; // @[G128Multiplay.scala 48:24:@3809.6]
  assign _T_1410 = _T_1406 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3815.6]
  assign V_63 = _T_1404 ? _T_1406 : _T_1410; // @[G128Multiplay.scala 46:7:@3808.4]
  assign _T_1412 = io_y[64]; // @[G128Multiplay.scala 37:16:@3819.4]
  assign _T_1415 = Z_63 ^ V_63; // @[G128Multiplay.scala 40:24:@3822.6]
  assign Z_64 = _T_1412 ? _T_1415 : Z_63; // @[G128Multiplay.scala 38:7:@3821.4]
  assign _T_1416 = V_63[0]; // @[G128Multiplay.scala 45:18:@3828.4]
  assign _T_1418 = _T_1416 == 1'h0; // @[G128Multiplay.scala 45:22:@3829.4]
  assign _T_1420 = V_63 >> 1'h1; // @[G128Multiplay.scala 48:24:@3831.6]
  assign _T_1424 = _T_1420 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3837.6]
  assign V_64 = _T_1418 ? _T_1420 : _T_1424; // @[G128Multiplay.scala 46:7:@3830.4]
  assign _T_1426 = io_y[63]; // @[G128Multiplay.scala 37:16:@3841.4]
  assign _T_1429 = Z_64 ^ V_64; // @[G128Multiplay.scala 40:24:@3844.6]
  assign Z_65 = _T_1426 ? _T_1429 : Z_64; // @[G128Multiplay.scala 38:7:@3843.4]
  assign _T_1430 = V_64[0]; // @[G128Multiplay.scala 45:18:@3850.4]
  assign _T_1432 = _T_1430 == 1'h0; // @[G128Multiplay.scala 45:22:@3851.4]
  assign _T_1434 = V_64 >> 1'h1; // @[G128Multiplay.scala 48:24:@3853.6]
  assign _T_1438 = _T_1434 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3859.6]
  assign V_65 = _T_1432 ? _T_1434 : _T_1438; // @[G128Multiplay.scala 46:7:@3852.4]
  assign _T_1440 = io_y[62]; // @[G128Multiplay.scala 37:16:@3863.4]
  assign _T_1443 = Z_65 ^ V_65; // @[G128Multiplay.scala 40:24:@3866.6]
  assign Z_66 = _T_1440 ? _T_1443 : Z_65; // @[G128Multiplay.scala 38:7:@3865.4]
  assign _T_1444 = V_65[0]; // @[G128Multiplay.scala 45:18:@3872.4]
  assign _T_1446 = _T_1444 == 1'h0; // @[G128Multiplay.scala 45:22:@3873.4]
  assign _T_1448 = V_65 >> 1'h1; // @[G128Multiplay.scala 48:24:@3875.6]
  assign _T_1452 = _T_1448 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3881.6]
  assign V_66 = _T_1446 ? _T_1448 : _T_1452; // @[G128Multiplay.scala 46:7:@3874.4]
  assign _T_1454 = io_y[61]; // @[G128Multiplay.scala 37:16:@3885.4]
  assign _T_1457 = Z_66 ^ V_66; // @[G128Multiplay.scala 40:24:@3888.6]
  assign Z_67 = _T_1454 ? _T_1457 : Z_66; // @[G128Multiplay.scala 38:7:@3887.4]
  assign _T_1458 = V_66[0]; // @[G128Multiplay.scala 45:18:@3894.4]
  assign _T_1460 = _T_1458 == 1'h0; // @[G128Multiplay.scala 45:22:@3895.4]
  assign _T_1462 = V_66 >> 1'h1; // @[G128Multiplay.scala 48:24:@3897.6]
  assign _T_1466 = _T_1462 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3903.6]
  assign V_67 = _T_1460 ? _T_1462 : _T_1466; // @[G128Multiplay.scala 46:7:@3896.4]
  assign _T_1468 = io_y[60]; // @[G128Multiplay.scala 37:16:@3907.4]
  assign _T_1471 = Z_67 ^ V_67; // @[G128Multiplay.scala 40:24:@3910.6]
  assign Z_68 = _T_1468 ? _T_1471 : Z_67; // @[G128Multiplay.scala 38:7:@3909.4]
  assign _T_1472 = V_67[0]; // @[G128Multiplay.scala 45:18:@3916.4]
  assign _T_1474 = _T_1472 == 1'h0; // @[G128Multiplay.scala 45:22:@3917.4]
  assign _T_1476 = V_67 >> 1'h1; // @[G128Multiplay.scala 48:24:@3919.6]
  assign _T_1480 = _T_1476 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3925.6]
  assign V_68 = _T_1474 ? _T_1476 : _T_1480; // @[G128Multiplay.scala 46:7:@3918.4]
  assign _T_1482 = io_y[59]; // @[G128Multiplay.scala 37:16:@3929.4]
  assign _T_1485 = Z_68 ^ V_68; // @[G128Multiplay.scala 40:24:@3932.6]
  assign Z_69 = _T_1482 ? _T_1485 : Z_68; // @[G128Multiplay.scala 38:7:@3931.4]
  assign _T_1486 = V_68[0]; // @[G128Multiplay.scala 45:18:@3938.4]
  assign _T_1488 = _T_1486 == 1'h0; // @[G128Multiplay.scala 45:22:@3939.4]
  assign _T_1490 = V_68 >> 1'h1; // @[G128Multiplay.scala 48:24:@3941.6]
  assign _T_1494 = _T_1490 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3947.6]
  assign V_69 = _T_1488 ? _T_1490 : _T_1494; // @[G128Multiplay.scala 46:7:@3940.4]
  assign _T_1496 = io_y[58]; // @[G128Multiplay.scala 37:16:@3951.4]
  assign _T_1499 = Z_69 ^ V_69; // @[G128Multiplay.scala 40:24:@3954.6]
  assign Z_70 = _T_1496 ? _T_1499 : Z_69; // @[G128Multiplay.scala 38:7:@3953.4]
  assign _T_1500 = V_69[0]; // @[G128Multiplay.scala 45:18:@3960.4]
  assign _T_1502 = _T_1500 == 1'h0; // @[G128Multiplay.scala 45:22:@3961.4]
  assign _T_1504 = V_69 >> 1'h1; // @[G128Multiplay.scala 48:24:@3963.6]
  assign _T_1508 = _T_1504 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3969.6]
  assign V_70 = _T_1502 ? _T_1504 : _T_1508; // @[G128Multiplay.scala 46:7:@3962.4]
  assign _T_1510 = io_y[57]; // @[G128Multiplay.scala 37:16:@3973.4]
  assign _T_1513 = Z_70 ^ V_70; // @[G128Multiplay.scala 40:24:@3976.6]
  assign Z_71 = _T_1510 ? _T_1513 : Z_70; // @[G128Multiplay.scala 38:7:@3975.4]
  assign _T_1514 = V_70[0]; // @[G128Multiplay.scala 45:18:@3982.4]
  assign _T_1516 = _T_1514 == 1'h0; // @[G128Multiplay.scala 45:22:@3983.4]
  assign _T_1518 = V_70 >> 1'h1; // @[G128Multiplay.scala 48:24:@3985.6]
  assign _T_1522 = _T_1518 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@3991.6]
  assign V_71 = _T_1516 ? _T_1518 : _T_1522; // @[G128Multiplay.scala 46:7:@3984.4]
  assign _T_1524 = io_y[56]; // @[G128Multiplay.scala 37:16:@3995.4]
  assign _T_1527 = Z_71 ^ V_71; // @[G128Multiplay.scala 40:24:@3998.6]
  assign Z_72 = _T_1524 ? _T_1527 : Z_71; // @[G128Multiplay.scala 38:7:@3997.4]
  assign _T_1528 = V_71[0]; // @[G128Multiplay.scala 45:18:@4004.4]
  assign _T_1530 = _T_1528 == 1'h0; // @[G128Multiplay.scala 45:22:@4005.4]
  assign _T_1532 = V_71 >> 1'h1; // @[G128Multiplay.scala 48:24:@4007.6]
  assign _T_1536 = _T_1532 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4013.6]
  assign V_72 = _T_1530 ? _T_1532 : _T_1536; // @[G128Multiplay.scala 46:7:@4006.4]
  assign _T_1538 = io_y[55]; // @[G128Multiplay.scala 37:16:@4017.4]
  assign _T_1541 = Z_72 ^ V_72; // @[G128Multiplay.scala 40:24:@4020.6]
  assign Z_73 = _T_1538 ? _T_1541 : Z_72; // @[G128Multiplay.scala 38:7:@4019.4]
  assign _T_1542 = V_72[0]; // @[G128Multiplay.scala 45:18:@4026.4]
  assign _T_1544 = _T_1542 == 1'h0; // @[G128Multiplay.scala 45:22:@4027.4]
  assign _T_1546 = V_72 >> 1'h1; // @[G128Multiplay.scala 48:24:@4029.6]
  assign _T_1550 = _T_1546 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4035.6]
  assign V_73 = _T_1544 ? _T_1546 : _T_1550; // @[G128Multiplay.scala 46:7:@4028.4]
  assign _T_1552 = io_y[54]; // @[G128Multiplay.scala 37:16:@4039.4]
  assign _T_1555 = Z_73 ^ V_73; // @[G128Multiplay.scala 40:24:@4042.6]
  assign Z_74 = _T_1552 ? _T_1555 : Z_73; // @[G128Multiplay.scala 38:7:@4041.4]
  assign _T_1556 = V_73[0]; // @[G128Multiplay.scala 45:18:@4048.4]
  assign _T_1558 = _T_1556 == 1'h0; // @[G128Multiplay.scala 45:22:@4049.4]
  assign _T_1560 = V_73 >> 1'h1; // @[G128Multiplay.scala 48:24:@4051.6]
  assign _T_1564 = _T_1560 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4057.6]
  assign V_74 = _T_1558 ? _T_1560 : _T_1564; // @[G128Multiplay.scala 46:7:@4050.4]
  assign _T_1566 = io_y[53]; // @[G128Multiplay.scala 37:16:@4061.4]
  assign _T_1569 = Z_74 ^ V_74; // @[G128Multiplay.scala 40:24:@4064.6]
  assign Z_75 = _T_1566 ? _T_1569 : Z_74; // @[G128Multiplay.scala 38:7:@4063.4]
  assign _T_1570 = V_74[0]; // @[G128Multiplay.scala 45:18:@4070.4]
  assign _T_1572 = _T_1570 == 1'h0; // @[G128Multiplay.scala 45:22:@4071.4]
  assign _T_1574 = V_74 >> 1'h1; // @[G128Multiplay.scala 48:24:@4073.6]
  assign _T_1578 = _T_1574 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4079.6]
  assign V_75 = _T_1572 ? _T_1574 : _T_1578; // @[G128Multiplay.scala 46:7:@4072.4]
  assign _T_1580 = io_y[52]; // @[G128Multiplay.scala 37:16:@4083.4]
  assign _T_1583 = Z_75 ^ V_75; // @[G128Multiplay.scala 40:24:@4086.6]
  assign Z_76 = _T_1580 ? _T_1583 : Z_75; // @[G128Multiplay.scala 38:7:@4085.4]
  assign _T_1584 = V_75[0]; // @[G128Multiplay.scala 45:18:@4092.4]
  assign _T_1586 = _T_1584 == 1'h0; // @[G128Multiplay.scala 45:22:@4093.4]
  assign _T_1588 = V_75 >> 1'h1; // @[G128Multiplay.scala 48:24:@4095.6]
  assign _T_1592 = _T_1588 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4101.6]
  assign V_76 = _T_1586 ? _T_1588 : _T_1592; // @[G128Multiplay.scala 46:7:@4094.4]
  assign _T_1594 = io_y[51]; // @[G128Multiplay.scala 37:16:@4105.4]
  assign _T_1597 = Z_76 ^ V_76; // @[G128Multiplay.scala 40:24:@4108.6]
  assign Z_77 = _T_1594 ? _T_1597 : Z_76; // @[G128Multiplay.scala 38:7:@4107.4]
  assign _T_1598 = V_76[0]; // @[G128Multiplay.scala 45:18:@4114.4]
  assign _T_1600 = _T_1598 == 1'h0; // @[G128Multiplay.scala 45:22:@4115.4]
  assign _T_1602 = V_76 >> 1'h1; // @[G128Multiplay.scala 48:24:@4117.6]
  assign _T_1606 = _T_1602 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4123.6]
  assign V_77 = _T_1600 ? _T_1602 : _T_1606; // @[G128Multiplay.scala 46:7:@4116.4]
  assign _T_1608 = io_y[50]; // @[G128Multiplay.scala 37:16:@4127.4]
  assign _T_1611 = Z_77 ^ V_77; // @[G128Multiplay.scala 40:24:@4130.6]
  assign Z_78 = _T_1608 ? _T_1611 : Z_77; // @[G128Multiplay.scala 38:7:@4129.4]
  assign _T_1612 = V_77[0]; // @[G128Multiplay.scala 45:18:@4136.4]
  assign _T_1614 = _T_1612 == 1'h0; // @[G128Multiplay.scala 45:22:@4137.4]
  assign _T_1616 = V_77 >> 1'h1; // @[G128Multiplay.scala 48:24:@4139.6]
  assign _T_1620 = _T_1616 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4145.6]
  assign V_78 = _T_1614 ? _T_1616 : _T_1620; // @[G128Multiplay.scala 46:7:@4138.4]
  assign _T_1622 = io_y[49]; // @[G128Multiplay.scala 37:16:@4149.4]
  assign _T_1625 = Z_78 ^ V_78; // @[G128Multiplay.scala 40:24:@4152.6]
  assign Z_79 = _T_1622 ? _T_1625 : Z_78; // @[G128Multiplay.scala 38:7:@4151.4]
  assign _T_1626 = V_78[0]; // @[G128Multiplay.scala 45:18:@4158.4]
  assign _T_1628 = _T_1626 == 1'h0; // @[G128Multiplay.scala 45:22:@4159.4]
  assign _T_1630 = V_78 >> 1'h1; // @[G128Multiplay.scala 48:24:@4161.6]
  assign _T_1634 = _T_1630 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4167.6]
  assign V_79 = _T_1628 ? _T_1630 : _T_1634; // @[G128Multiplay.scala 46:7:@4160.4]
  assign _T_1636 = io_y[48]; // @[G128Multiplay.scala 37:16:@4171.4]
  assign _T_1639 = Z_79 ^ V_79; // @[G128Multiplay.scala 40:24:@4174.6]
  assign Z_80 = _T_1636 ? _T_1639 : Z_79; // @[G128Multiplay.scala 38:7:@4173.4]
  assign _T_1640 = V_79[0]; // @[G128Multiplay.scala 45:18:@4180.4]
  assign _T_1642 = _T_1640 == 1'h0; // @[G128Multiplay.scala 45:22:@4181.4]
  assign _T_1644 = V_79 >> 1'h1; // @[G128Multiplay.scala 48:24:@4183.6]
  assign _T_1648 = _T_1644 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4189.6]
  assign V_80 = _T_1642 ? _T_1644 : _T_1648; // @[G128Multiplay.scala 46:7:@4182.4]
  assign _T_1650 = io_y[47]; // @[G128Multiplay.scala 37:16:@4193.4]
  assign _T_1653 = Z_80 ^ V_80; // @[G128Multiplay.scala 40:24:@4196.6]
  assign Z_81 = _T_1650 ? _T_1653 : Z_80; // @[G128Multiplay.scala 38:7:@4195.4]
  assign _T_1654 = V_80[0]; // @[G128Multiplay.scala 45:18:@4202.4]
  assign _T_1656 = _T_1654 == 1'h0; // @[G128Multiplay.scala 45:22:@4203.4]
  assign _T_1658 = V_80 >> 1'h1; // @[G128Multiplay.scala 48:24:@4205.6]
  assign _T_1662 = _T_1658 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4211.6]
  assign V_81 = _T_1656 ? _T_1658 : _T_1662; // @[G128Multiplay.scala 46:7:@4204.4]
  assign _T_1664 = io_y[46]; // @[G128Multiplay.scala 37:16:@4215.4]
  assign _T_1667 = Z_81 ^ V_81; // @[G128Multiplay.scala 40:24:@4218.6]
  assign Z_82 = _T_1664 ? _T_1667 : Z_81; // @[G128Multiplay.scala 38:7:@4217.4]
  assign _T_1668 = V_81[0]; // @[G128Multiplay.scala 45:18:@4224.4]
  assign _T_1670 = _T_1668 == 1'h0; // @[G128Multiplay.scala 45:22:@4225.4]
  assign _T_1672 = V_81 >> 1'h1; // @[G128Multiplay.scala 48:24:@4227.6]
  assign _T_1676 = _T_1672 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4233.6]
  assign V_82 = _T_1670 ? _T_1672 : _T_1676; // @[G128Multiplay.scala 46:7:@4226.4]
  assign _T_1678 = io_y[45]; // @[G128Multiplay.scala 37:16:@4237.4]
  assign _T_1681 = Z_82 ^ V_82; // @[G128Multiplay.scala 40:24:@4240.6]
  assign Z_83 = _T_1678 ? _T_1681 : Z_82; // @[G128Multiplay.scala 38:7:@4239.4]
  assign _T_1682 = V_82[0]; // @[G128Multiplay.scala 45:18:@4246.4]
  assign _T_1684 = _T_1682 == 1'h0; // @[G128Multiplay.scala 45:22:@4247.4]
  assign _T_1686 = V_82 >> 1'h1; // @[G128Multiplay.scala 48:24:@4249.6]
  assign _T_1690 = _T_1686 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4255.6]
  assign V_83 = _T_1684 ? _T_1686 : _T_1690; // @[G128Multiplay.scala 46:7:@4248.4]
  assign _T_1692 = io_y[44]; // @[G128Multiplay.scala 37:16:@4259.4]
  assign _T_1695 = Z_83 ^ V_83; // @[G128Multiplay.scala 40:24:@4262.6]
  assign Z_84 = _T_1692 ? _T_1695 : Z_83; // @[G128Multiplay.scala 38:7:@4261.4]
  assign _T_1696 = V_83[0]; // @[G128Multiplay.scala 45:18:@4268.4]
  assign _T_1698 = _T_1696 == 1'h0; // @[G128Multiplay.scala 45:22:@4269.4]
  assign _T_1700 = V_83 >> 1'h1; // @[G128Multiplay.scala 48:24:@4271.6]
  assign _T_1704 = _T_1700 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4277.6]
  assign V_84 = _T_1698 ? _T_1700 : _T_1704; // @[G128Multiplay.scala 46:7:@4270.4]
  assign _T_1706 = io_y[43]; // @[G128Multiplay.scala 37:16:@4281.4]
  assign _T_1709 = Z_84 ^ V_84; // @[G128Multiplay.scala 40:24:@4284.6]
  assign Z_85 = _T_1706 ? _T_1709 : Z_84; // @[G128Multiplay.scala 38:7:@4283.4]
  assign _T_1710 = V_84[0]; // @[G128Multiplay.scala 45:18:@4290.4]
  assign _T_1712 = _T_1710 == 1'h0; // @[G128Multiplay.scala 45:22:@4291.4]
  assign _T_1714 = V_84 >> 1'h1; // @[G128Multiplay.scala 48:24:@4293.6]
  assign _T_1718 = _T_1714 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4299.6]
  assign V_85 = _T_1712 ? _T_1714 : _T_1718; // @[G128Multiplay.scala 46:7:@4292.4]
  assign _T_1720 = io_y[42]; // @[G128Multiplay.scala 37:16:@4303.4]
  assign _T_1723 = Z_85 ^ V_85; // @[G128Multiplay.scala 40:24:@4306.6]
  assign Z_86 = _T_1720 ? _T_1723 : Z_85; // @[G128Multiplay.scala 38:7:@4305.4]
  assign _T_1724 = V_85[0]; // @[G128Multiplay.scala 45:18:@4312.4]
  assign _T_1726 = _T_1724 == 1'h0; // @[G128Multiplay.scala 45:22:@4313.4]
  assign _T_1728 = V_85 >> 1'h1; // @[G128Multiplay.scala 48:24:@4315.6]
  assign _T_1732 = _T_1728 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4321.6]
  assign V_86 = _T_1726 ? _T_1728 : _T_1732; // @[G128Multiplay.scala 46:7:@4314.4]
  assign _T_1734 = io_y[41]; // @[G128Multiplay.scala 37:16:@4325.4]
  assign _T_1737 = Z_86 ^ V_86; // @[G128Multiplay.scala 40:24:@4328.6]
  assign Z_87 = _T_1734 ? _T_1737 : Z_86; // @[G128Multiplay.scala 38:7:@4327.4]
  assign _T_1738 = V_86[0]; // @[G128Multiplay.scala 45:18:@4334.4]
  assign _T_1740 = _T_1738 == 1'h0; // @[G128Multiplay.scala 45:22:@4335.4]
  assign _T_1742 = V_86 >> 1'h1; // @[G128Multiplay.scala 48:24:@4337.6]
  assign _T_1746 = _T_1742 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4343.6]
  assign V_87 = _T_1740 ? _T_1742 : _T_1746; // @[G128Multiplay.scala 46:7:@4336.4]
  assign _T_1748 = io_y[40]; // @[G128Multiplay.scala 37:16:@4347.4]
  assign _T_1751 = Z_87 ^ V_87; // @[G128Multiplay.scala 40:24:@4350.6]
  assign Z_88 = _T_1748 ? _T_1751 : Z_87; // @[G128Multiplay.scala 38:7:@4349.4]
  assign _T_1752 = V_87[0]; // @[G128Multiplay.scala 45:18:@4356.4]
  assign _T_1754 = _T_1752 == 1'h0; // @[G128Multiplay.scala 45:22:@4357.4]
  assign _T_1756 = V_87 >> 1'h1; // @[G128Multiplay.scala 48:24:@4359.6]
  assign _T_1760 = _T_1756 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4365.6]
  assign V_88 = _T_1754 ? _T_1756 : _T_1760; // @[G128Multiplay.scala 46:7:@4358.4]
  assign _T_1762 = io_y[39]; // @[G128Multiplay.scala 37:16:@4369.4]
  assign _T_1765 = Z_88 ^ V_88; // @[G128Multiplay.scala 40:24:@4372.6]
  assign Z_89 = _T_1762 ? _T_1765 : Z_88; // @[G128Multiplay.scala 38:7:@4371.4]
  assign _T_1766 = V_88[0]; // @[G128Multiplay.scala 45:18:@4378.4]
  assign _T_1768 = _T_1766 == 1'h0; // @[G128Multiplay.scala 45:22:@4379.4]
  assign _T_1770 = V_88 >> 1'h1; // @[G128Multiplay.scala 48:24:@4381.6]
  assign _T_1774 = _T_1770 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4387.6]
  assign V_89 = _T_1768 ? _T_1770 : _T_1774; // @[G128Multiplay.scala 46:7:@4380.4]
  assign _T_1776 = io_y[38]; // @[G128Multiplay.scala 37:16:@4391.4]
  assign _T_1779 = Z_89 ^ V_89; // @[G128Multiplay.scala 40:24:@4394.6]
  assign Z_90 = _T_1776 ? _T_1779 : Z_89; // @[G128Multiplay.scala 38:7:@4393.4]
  assign _T_1780 = V_89[0]; // @[G128Multiplay.scala 45:18:@4400.4]
  assign _T_1782 = _T_1780 == 1'h0; // @[G128Multiplay.scala 45:22:@4401.4]
  assign _T_1784 = V_89 >> 1'h1; // @[G128Multiplay.scala 48:24:@4403.6]
  assign _T_1788 = _T_1784 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4409.6]
  assign V_90 = _T_1782 ? _T_1784 : _T_1788; // @[G128Multiplay.scala 46:7:@4402.4]
  assign _T_1790 = io_y[37]; // @[G128Multiplay.scala 37:16:@4413.4]
  assign _T_1793 = Z_90 ^ V_90; // @[G128Multiplay.scala 40:24:@4416.6]
  assign Z_91 = _T_1790 ? _T_1793 : Z_90; // @[G128Multiplay.scala 38:7:@4415.4]
  assign _T_1794 = V_90[0]; // @[G128Multiplay.scala 45:18:@4422.4]
  assign _T_1796 = _T_1794 == 1'h0; // @[G128Multiplay.scala 45:22:@4423.4]
  assign _T_1798 = V_90 >> 1'h1; // @[G128Multiplay.scala 48:24:@4425.6]
  assign _T_1802 = _T_1798 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4431.6]
  assign V_91 = _T_1796 ? _T_1798 : _T_1802; // @[G128Multiplay.scala 46:7:@4424.4]
  assign _T_1804 = io_y[36]; // @[G128Multiplay.scala 37:16:@4435.4]
  assign _T_1807 = Z_91 ^ V_91; // @[G128Multiplay.scala 40:24:@4438.6]
  assign Z_92 = _T_1804 ? _T_1807 : Z_91; // @[G128Multiplay.scala 38:7:@4437.4]
  assign _T_1808 = V_91[0]; // @[G128Multiplay.scala 45:18:@4444.4]
  assign _T_1810 = _T_1808 == 1'h0; // @[G128Multiplay.scala 45:22:@4445.4]
  assign _T_1812 = V_91 >> 1'h1; // @[G128Multiplay.scala 48:24:@4447.6]
  assign _T_1816 = _T_1812 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4453.6]
  assign V_92 = _T_1810 ? _T_1812 : _T_1816; // @[G128Multiplay.scala 46:7:@4446.4]
  assign _T_1818 = io_y[35]; // @[G128Multiplay.scala 37:16:@4457.4]
  assign _T_1821 = Z_92 ^ V_92; // @[G128Multiplay.scala 40:24:@4460.6]
  assign Z_93 = _T_1818 ? _T_1821 : Z_92; // @[G128Multiplay.scala 38:7:@4459.4]
  assign _T_1822 = V_92[0]; // @[G128Multiplay.scala 45:18:@4466.4]
  assign _T_1824 = _T_1822 == 1'h0; // @[G128Multiplay.scala 45:22:@4467.4]
  assign _T_1826 = V_92 >> 1'h1; // @[G128Multiplay.scala 48:24:@4469.6]
  assign _T_1830 = _T_1826 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4475.6]
  assign V_93 = _T_1824 ? _T_1826 : _T_1830; // @[G128Multiplay.scala 46:7:@4468.4]
  assign _T_1832 = io_y[34]; // @[G128Multiplay.scala 37:16:@4479.4]
  assign _T_1835 = Z_93 ^ V_93; // @[G128Multiplay.scala 40:24:@4482.6]
  assign Z_94 = _T_1832 ? _T_1835 : Z_93; // @[G128Multiplay.scala 38:7:@4481.4]
  assign _T_1836 = V_93[0]; // @[G128Multiplay.scala 45:18:@4488.4]
  assign _T_1838 = _T_1836 == 1'h0; // @[G128Multiplay.scala 45:22:@4489.4]
  assign _T_1840 = V_93 >> 1'h1; // @[G128Multiplay.scala 48:24:@4491.6]
  assign _T_1844 = _T_1840 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4497.6]
  assign V_94 = _T_1838 ? _T_1840 : _T_1844; // @[G128Multiplay.scala 46:7:@4490.4]
  assign _T_1846 = io_y[33]; // @[G128Multiplay.scala 37:16:@4501.4]
  assign _T_1849 = Z_94 ^ V_94; // @[G128Multiplay.scala 40:24:@4504.6]
  assign Z_95 = _T_1846 ? _T_1849 : Z_94; // @[G128Multiplay.scala 38:7:@4503.4]
  assign _T_1850 = V_94[0]; // @[G128Multiplay.scala 45:18:@4510.4]
  assign _T_1852 = _T_1850 == 1'h0; // @[G128Multiplay.scala 45:22:@4511.4]
  assign _T_1854 = V_94 >> 1'h1; // @[G128Multiplay.scala 48:24:@4513.6]
  assign _T_1858 = _T_1854 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4519.6]
  assign V_95 = _T_1852 ? _T_1854 : _T_1858; // @[G128Multiplay.scala 46:7:@4512.4]
  assign _T_1860 = io_y[32]; // @[G128Multiplay.scala 37:16:@4523.4]
  assign _T_1863 = Z_95 ^ V_95; // @[G128Multiplay.scala 40:24:@4526.6]
  assign Z_96 = _T_1860 ? _T_1863 : Z_95; // @[G128Multiplay.scala 38:7:@4525.4]
  assign _T_1864 = V_95[0]; // @[G128Multiplay.scala 45:18:@4532.4]
  assign _T_1866 = _T_1864 == 1'h0; // @[G128Multiplay.scala 45:22:@4533.4]
  assign _T_1868 = V_95 >> 1'h1; // @[G128Multiplay.scala 48:24:@4535.6]
  assign _T_1872 = _T_1868 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4541.6]
  assign V_96 = _T_1866 ? _T_1868 : _T_1872; // @[G128Multiplay.scala 46:7:@4534.4]
  assign _T_1874 = io_y[31]; // @[G128Multiplay.scala 37:16:@4545.4]
  assign _T_1877 = Z_96 ^ V_96; // @[G128Multiplay.scala 40:24:@4548.6]
  assign Z_97 = _T_1874 ? _T_1877 : Z_96; // @[G128Multiplay.scala 38:7:@4547.4]
  assign _T_1878 = V_96[0]; // @[G128Multiplay.scala 45:18:@4554.4]
  assign _T_1880 = _T_1878 == 1'h0; // @[G128Multiplay.scala 45:22:@4555.4]
  assign _T_1882 = V_96 >> 1'h1; // @[G128Multiplay.scala 48:24:@4557.6]
  assign _T_1886 = _T_1882 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4563.6]
  assign V_97 = _T_1880 ? _T_1882 : _T_1886; // @[G128Multiplay.scala 46:7:@4556.4]
  assign _T_1888 = io_y[30]; // @[G128Multiplay.scala 37:16:@4567.4]
  assign _T_1891 = Z_97 ^ V_97; // @[G128Multiplay.scala 40:24:@4570.6]
  assign Z_98 = _T_1888 ? _T_1891 : Z_97; // @[G128Multiplay.scala 38:7:@4569.4]
  assign _T_1892 = V_97[0]; // @[G128Multiplay.scala 45:18:@4576.4]
  assign _T_1894 = _T_1892 == 1'h0; // @[G128Multiplay.scala 45:22:@4577.4]
  assign _T_1896 = V_97 >> 1'h1; // @[G128Multiplay.scala 48:24:@4579.6]
  assign _T_1900 = _T_1896 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4585.6]
  assign V_98 = _T_1894 ? _T_1896 : _T_1900; // @[G128Multiplay.scala 46:7:@4578.4]
  assign _T_1902 = io_y[29]; // @[G128Multiplay.scala 37:16:@4589.4]
  assign _T_1905 = Z_98 ^ V_98; // @[G128Multiplay.scala 40:24:@4592.6]
  assign Z_99 = _T_1902 ? _T_1905 : Z_98; // @[G128Multiplay.scala 38:7:@4591.4]
  assign _T_1906 = V_98[0]; // @[G128Multiplay.scala 45:18:@4598.4]
  assign _T_1908 = _T_1906 == 1'h0; // @[G128Multiplay.scala 45:22:@4599.4]
  assign _T_1910 = V_98 >> 1'h1; // @[G128Multiplay.scala 48:24:@4601.6]
  assign _T_1914 = _T_1910 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4607.6]
  assign V_99 = _T_1908 ? _T_1910 : _T_1914; // @[G128Multiplay.scala 46:7:@4600.4]
  assign _T_1916 = io_y[28]; // @[G128Multiplay.scala 37:16:@4611.4]
  assign _T_1919 = Z_99 ^ V_99; // @[G128Multiplay.scala 40:24:@4614.6]
  assign Z_100 = _T_1916 ? _T_1919 : Z_99; // @[G128Multiplay.scala 38:7:@4613.4]
  assign _T_1920 = V_99[0]; // @[G128Multiplay.scala 45:18:@4620.4]
  assign _T_1922 = _T_1920 == 1'h0; // @[G128Multiplay.scala 45:22:@4621.4]
  assign _T_1924 = V_99 >> 1'h1; // @[G128Multiplay.scala 48:24:@4623.6]
  assign _T_1928 = _T_1924 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4629.6]
  assign V_100 = _T_1922 ? _T_1924 : _T_1928; // @[G128Multiplay.scala 46:7:@4622.4]
  assign _T_1930 = io_y[27]; // @[G128Multiplay.scala 37:16:@4633.4]
  assign _T_1933 = Z_100 ^ V_100; // @[G128Multiplay.scala 40:24:@4636.6]
  assign Z_101 = _T_1930 ? _T_1933 : Z_100; // @[G128Multiplay.scala 38:7:@4635.4]
  assign _T_1934 = V_100[0]; // @[G128Multiplay.scala 45:18:@4642.4]
  assign _T_1936 = _T_1934 == 1'h0; // @[G128Multiplay.scala 45:22:@4643.4]
  assign _T_1938 = V_100 >> 1'h1; // @[G128Multiplay.scala 48:24:@4645.6]
  assign _T_1942 = _T_1938 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4651.6]
  assign V_101 = _T_1936 ? _T_1938 : _T_1942; // @[G128Multiplay.scala 46:7:@4644.4]
  assign _T_1944 = io_y[26]; // @[G128Multiplay.scala 37:16:@4655.4]
  assign _T_1947 = Z_101 ^ V_101; // @[G128Multiplay.scala 40:24:@4658.6]
  assign Z_102 = _T_1944 ? _T_1947 : Z_101; // @[G128Multiplay.scala 38:7:@4657.4]
  assign _T_1948 = V_101[0]; // @[G128Multiplay.scala 45:18:@4664.4]
  assign _T_1950 = _T_1948 == 1'h0; // @[G128Multiplay.scala 45:22:@4665.4]
  assign _T_1952 = V_101 >> 1'h1; // @[G128Multiplay.scala 48:24:@4667.6]
  assign _T_1956 = _T_1952 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4673.6]
  assign V_102 = _T_1950 ? _T_1952 : _T_1956; // @[G128Multiplay.scala 46:7:@4666.4]
  assign _T_1958 = io_y[25]; // @[G128Multiplay.scala 37:16:@4677.4]
  assign _T_1961 = Z_102 ^ V_102; // @[G128Multiplay.scala 40:24:@4680.6]
  assign Z_103 = _T_1958 ? _T_1961 : Z_102; // @[G128Multiplay.scala 38:7:@4679.4]
  assign _T_1962 = V_102[0]; // @[G128Multiplay.scala 45:18:@4686.4]
  assign _T_1964 = _T_1962 == 1'h0; // @[G128Multiplay.scala 45:22:@4687.4]
  assign _T_1966 = V_102 >> 1'h1; // @[G128Multiplay.scala 48:24:@4689.6]
  assign _T_1970 = _T_1966 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4695.6]
  assign V_103 = _T_1964 ? _T_1966 : _T_1970; // @[G128Multiplay.scala 46:7:@4688.4]
  assign _T_1972 = io_y[24]; // @[G128Multiplay.scala 37:16:@4699.4]
  assign _T_1975 = Z_103 ^ V_103; // @[G128Multiplay.scala 40:24:@4702.6]
  assign Z_104 = _T_1972 ? _T_1975 : Z_103; // @[G128Multiplay.scala 38:7:@4701.4]
  assign _T_1976 = V_103[0]; // @[G128Multiplay.scala 45:18:@4708.4]
  assign _T_1978 = _T_1976 == 1'h0; // @[G128Multiplay.scala 45:22:@4709.4]
  assign _T_1980 = V_103 >> 1'h1; // @[G128Multiplay.scala 48:24:@4711.6]
  assign _T_1984 = _T_1980 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4717.6]
  assign V_104 = _T_1978 ? _T_1980 : _T_1984; // @[G128Multiplay.scala 46:7:@4710.4]
  assign _T_1986 = io_y[23]; // @[G128Multiplay.scala 37:16:@4721.4]
  assign _T_1989 = Z_104 ^ V_104; // @[G128Multiplay.scala 40:24:@4724.6]
  assign Z_105 = _T_1986 ? _T_1989 : Z_104; // @[G128Multiplay.scala 38:7:@4723.4]
  assign _T_1990 = V_104[0]; // @[G128Multiplay.scala 45:18:@4730.4]
  assign _T_1992 = _T_1990 == 1'h0; // @[G128Multiplay.scala 45:22:@4731.4]
  assign _T_1994 = V_104 >> 1'h1; // @[G128Multiplay.scala 48:24:@4733.6]
  assign _T_1998 = _T_1994 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4739.6]
  assign V_105 = _T_1992 ? _T_1994 : _T_1998; // @[G128Multiplay.scala 46:7:@4732.4]
  assign _T_2000 = io_y[22]; // @[G128Multiplay.scala 37:16:@4743.4]
  assign _T_2003 = Z_105 ^ V_105; // @[G128Multiplay.scala 40:24:@4746.6]
  assign Z_106 = _T_2000 ? _T_2003 : Z_105; // @[G128Multiplay.scala 38:7:@4745.4]
  assign _T_2004 = V_105[0]; // @[G128Multiplay.scala 45:18:@4752.4]
  assign _T_2006 = _T_2004 == 1'h0; // @[G128Multiplay.scala 45:22:@4753.4]
  assign _T_2008 = V_105 >> 1'h1; // @[G128Multiplay.scala 48:24:@4755.6]
  assign _T_2012 = _T_2008 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4761.6]
  assign V_106 = _T_2006 ? _T_2008 : _T_2012; // @[G128Multiplay.scala 46:7:@4754.4]
  assign _T_2014 = io_y[21]; // @[G128Multiplay.scala 37:16:@4765.4]
  assign _T_2017 = Z_106 ^ V_106; // @[G128Multiplay.scala 40:24:@4768.6]
  assign Z_107 = _T_2014 ? _T_2017 : Z_106; // @[G128Multiplay.scala 38:7:@4767.4]
  assign _T_2018 = V_106[0]; // @[G128Multiplay.scala 45:18:@4774.4]
  assign _T_2020 = _T_2018 == 1'h0; // @[G128Multiplay.scala 45:22:@4775.4]
  assign _T_2022 = V_106 >> 1'h1; // @[G128Multiplay.scala 48:24:@4777.6]
  assign _T_2026 = _T_2022 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4783.6]
  assign V_107 = _T_2020 ? _T_2022 : _T_2026; // @[G128Multiplay.scala 46:7:@4776.4]
  assign _T_2028 = io_y[20]; // @[G128Multiplay.scala 37:16:@4787.4]
  assign _T_2031 = Z_107 ^ V_107; // @[G128Multiplay.scala 40:24:@4790.6]
  assign Z_108 = _T_2028 ? _T_2031 : Z_107; // @[G128Multiplay.scala 38:7:@4789.4]
  assign _T_2032 = V_107[0]; // @[G128Multiplay.scala 45:18:@4796.4]
  assign _T_2034 = _T_2032 == 1'h0; // @[G128Multiplay.scala 45:22:@4797.4]
  assign _T_2036 = V_107 >> 1'h1; // @[G128Multiplay.scala 48:24:@4799.6]
  assign _T_2040 = _T_2036 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4805.6]
  assign V_108 = _T_2034 ? _T_2036 : _T_2040; // @[G128Multiplay.scala 46:7:@4798.4]
  assign _T_2042 = io_y[19]; // @[G128Multiplay.scala 37:16:@4809.4]
  assign _T_2045 = Z_108 ^ V_108; // @[G128Multiplay.scala 40:24:@4812.6]
  assign Z_109 = _T_2042 ? _T_2045 : Z_108; // @[G128Multiplay.scala 38:7:@4811.4]
  assign _T_2046 = V_108[0]; // @[G128Multiplay.scala 45:18:@4818.4]
  assign _T_2048 = _T_2046 == 1'h0; // @[G128Multiplay.scala 45:22:@4819.4]
  assign _T_2050 = V_108 >> 1'h1; // @[G128Multiplay.scala 48:24:@4821.6]
  assign _T_2054 = _T_2050 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4827.6]
  assign V_109 = _T_2048 ? _T_2050 : _T_2054; // @[G128Multiplay.scala 46:7:@4820.4]
  assign _T_2056 = io_y[18]; // @[G128Multiplay.scala 37:16:@4831.4]
  assign _T_2059 = Z_109 ^ V_109; // @[G128Multiplay.scala 40:24:@4834.6]
  assign Z_110 = _T_2056 ? _T_2059 : Z_109; // @[G128Multiplay.scala 38:7:@4833.4]
  assign _T_2060 = V_109[0]; // @[G128Multiplay.scala 45:18:@4840.4]
  assign _T_2062 = _T_2060 == 1'h0; // @[G128Multiplay.scala 45:22:@4841.4]
  assign _T_2064 = V_109 >> 1'h1; // @[G128Multiplay.scala 48:24:@4843.6]
  assign _T_2068 = _T_2064 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4849.6]
  assign V_110 = _T_2062 ? _T_2064 : _T_2068; // @[G128Multiplay.scala 46:7:@4842.4]
  assign _T_2070 = io_y[17]; // @[G128Multiplay.scala 37:16:@4853.4]
  assign _T_2073 = Z_110 ^ V_110; // @[G128Multiplay.scala 40:24:@4856.6]
  assign Z_111 = _T_2070 ? _T_2073 : Z_110; // @[G128Multiplay.scala 38:7:@4855.4]
  assign _T_2074 = V_110[0]; // @[G128Multiplay.scala 45:18:@4862.4]
  assign _T_2076 = _T_2074 == 1'h0; // @[G128Multiplay.scala 45:22:@4863.4]
  assign _T_2078 = V_110 >> 1'h1; // @[G128Multiplay.scala 48:24:@4865.6]
  assign _T_2082 = _T_2078 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4871.6]
  assign V_111 = _T_2076 ? _T_2078 : _T_2082; // @[G128Multiplay.scala 46:7:@4864.4]
  assign _T_2084 = io_y[16]; // @[G128Multiplay.scala 37:16:@4875.4]
  assign _T_2087 = Z_111 ^ V_111; // @[G128Multiplay.scala 40:24:@4878.6]
  assign Z_112 = _T_2084 ? _T_2087 : Z_111; // @[G128Multiplay.scala 38:7:@4877.4]
  assign _T_2088 = V_111[0]; // @[G128Multiplay.scala 45:18:@4884.4]
  assign _T_2090 = _T_2088 == 1'h0; // @[G128Multiplay.scala 45:22:@4885.4]
  assign _T_2092 = V_111 >> 1'h1; // @[G128Multiplay.scala 48:24:@4887.6]
  assign _T_2096 = _T_2092 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4893.6]
  assign V_112 = _T_2090 ? _T_2092 : _T_2096; // @[G128Multiplay.scala 46:7:@4886.4]
  assign _T_2098 = io_y[15]; // @[G128Multiplay.scala 37:16:@4897.4]
  assign _T_2101 = Z_112 ^ V_112; // @[G128Multiplay.scala 40:24:@4900.6]
  assign Z_113 = _T_2098 ? _T_2101 : Z_112; // @[G128Multiplay.scala 38:7:@4899.4]
  assign _T_2102 = V_112[0]; // @[G128Multiplay.scala 45:18:@4906.4]
  assign _T_2104 = _T_2102 == 1'h0; // @[G128Multiplay.scala 45:22:@4907.4]
  assign _T_2106 = V_112 >> 1'h1; // @[G128Multiplay.scala 48:24:@4909.6]
  assign _T_2110 = _T_2106 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4915.6]
  assign V_113 = _T_2104 ? _T_2106 : _T_2110; // @[G128Multiplay.scala 46:7:@4908.4]
  assign _T_2112 = io_y[14]; // @[G128Multiplay.scala 37:16:@4919.4]
  assign _T_2115 = Z_113 ^ V_113; // @[G128Multiplay.scala 40:24:@4922.6]
  assign Z_114 = _T_2112 ? _T_2115 : Z_113; // @[G128Multiplay.scala 38:7:@4921.4]
  assign _T_2116 = V_113[0]; // @[G128Multiplay.scala 45:18:@4928.4]
  assign _T_2118 = _T_2116 == 1'h0; // @[G128Multiplay.scala 45:22:@4929.4]
  assign _T_2120 = V_113 >> 1'h1; // @[G128Multiplay.scala 48:24:@4931.6]
  assign _T_2124 = _T_2120 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4937.6]
  assign V_114 = _T_2118 ? _T_2120 : _T_2124; // @[G128Multiplay.scala 46:7:@4930.4]
  assign _T_2126 = io_y[13]; // @[G128Multiplay.scala 37:16:@4941.4]
  assign _T_2129 = Z_114 ^ V_114; // @[G128Multiplay.scala 40:24:@4944.6]
  assign Z_115 = _T_2126 ? _T_2129 : Z_114; // @[G128Multiplay.scala 38:7:@4943.4]
  assign _T_2130 = V_114[0]; // @[G128Multiplay.scala 45:18:@4950.4]
  assign _T_2132 = _T_2130 == 1'h0; // @[G128Multiplay.scala 45:22:@4951.4]
  assign _T_2134 = V_114 >> 1'h1; // @[G128Multiplay.scala 48:24:@4953.6]
  assign _T_2138 = _T_2134 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4959.6]
  assign V_115 = _T_2132 ? _T_2134 : _T_2138; // @[G128Multiplay.scala 46:7:@4952.4]
  assign _T_2140 = io_y[12]; // @[G128Multiplay.scala 37:16:@4963.4]
  assign _T_2143 = Z_115 ^ V_115; // @[G128Multiplay.scala 40:24:@4966.6]
  assign Z_116 = _T_2140 ? _T_2143 : Z_115; // @[G128Multiplay.scala 38:7:@4965.4]
  assign _T_2144 = V_115[0]; // @[G128Multiplay.scala 45:18:@4972.4]
  assign _T_2146 = _T_2144 == 1'h0; // @[G128Multiplay.scala 45:22:@4973.4]
  assign _T_2148 = V_115 >> 1'h1; // @[G128Multiplay.scala 48:24:@4975.6]
  assign _T_2152 = _T_2148 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@4981.6]
  assign V_116 = _T_2146 ? _T_2148 : _T_2152; // @[G128Multiplay.scala 46:7:@4974.4]
  assign _T_2154 = io_y[11]; // @[G128Multiplay.scala 37:16:@4985.4]
  assign _T_2157 = Z_116 ^ V_116; // @[G128Multiplay.scala 40:24:@4988.6]
  assign Z_117 = _T_2154 ? _T_2157 : Z_116; // @[G128Multiplay.scala 38:7:@4987.4]
  assign _T_2158 = V_116[0]; // @[G128Multiplay.scala 45:18:@4994.4]
  assign _T_2160 = _T_2158 == 1'h0; // @[G128Multiplay.scala 45:22:@4995.4]
  assign _T_2162 = V_116 >> 1'h1; // @[G128Multiplay.scala 48:24:@4997.6]
  assign _T_2166 = _T_2162 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5003.6]
  assign V_117 = _T_2160 ? _T_2162 : _T_2166; // @[G128Multiplay.scala 46:7:@4996.4]
  assign _T_2168 = io_y[10]; // @[G128Multiplay.scala 37:16:@5007.4]
  assign _T_2171 = Z_117 ^ V_117; // @[G128Multiplay.scala 40:24:@5010.6]
  assign Z_118 = _T_2168 ? _T_2171 : Z_117; // @[G128Multiplay.scala 38:7:@5009.4]
  assign _T_2172 = V_117[0]; // @[G128Multiplay.scala 45:18:@5016.4]
  assign _T_2174 = _T_2172 == 1'h0; // @[G128Multiplay.scala 45:22:@5017.4]
  assign _T_2176 = V_117 >> 1'h1; // @[G128Multiplay.scala 48:24:@5019.6]
  assign _T_2180 = _T_2176 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5025.6]
  assign V_118 = _T_2174 ? _T_2176 : _T_2180; // @[G128Multiplay.scala 46:7:@5018.4]
  assign _T_2182 = io_y[9]; // @[G128Multiplay.scala 37:16:@5029.4]
  assign _T_2185 = Z_118 ^ V_118; // @[G128Multiplay.scala 40:24:@5032.6]
  assign Z_119 = _T_2182 ? _T_2185 : Z_118; // @[G128Multiplay.scala 38:7:@5031.4]
  assign _T_2186 = V_118[0]; // @[G128Multiplay.scala 45:18:@5038.4]
  assign _T_2188 = _T_2186 == 1'h0; // @[G128Multiplay.scala 45:22:@5039.4]
  assign _T_2190 = V_118 >> 1'h1; // @[G128Multiplay.scala 48:24:@5041.6]
  assign _T_2194 = _T_2190 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5047.6]
  assign V_119 = _T_2188 ? _T_2190 : _T_2194; // @[G128Multiplay.scala 46:7:@5040.4]
  assign _T_2196 = io_y[8]; // @[G128Multiplay.scala 37:16:@5051.4]
  assign _T_2199 = Z_119 ^ V_119; // @[G128Multiplay.scala 40:24:@5054.6]
  assign Z_120 = _T_2196 ? _T_2199 : Z_119; // @[G128Multiplay.scala 38:7:@5053.4]
  assign _T_2200 = V_119[0]; // @[G128Multiplay.scala 45:18:@5060.4]
  assign _T_2202 = _T_2200 == 1'h0; // @[G128Multiplay.scala 45:22:@5061.4]
  assign _T_2204 = V_119 >> 1'h1; // @[G128Multiplay.scala 48:24:@5063.6]
  assign _T_2208 = _T_2204 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5069.6]
  assign V_120 = _T_2202 ? _T_2204 : _T_2208; // @[G128Multiplay.scala 46:7:@5062.4]
  assign _T_2210 = io_y[7]; // @[G128Multiplay.scala 37:16:@5073.4]
  assign _T_2213 = Z_120 ^ V_120; // @[G128Multiplay.scala 40:24:@5076.6]
  assign Z_121 = _T_2210 ? _T_2213 : Z_120; // @[G128Multiplay.scala 38:7:@5075.4]
  assign _T_2214 = V_120[0]; // @[G128Multiplay.scala 45:18:@5082.4]
  assign _T_2216 = _T_2214 == 1'h0; // @[G128Multiplay.scala 45:22:@5083.4]
  assign _T_2218 = V_120 >> 1'h1; // @[G128Multiplay.scala 48:24:@5085.6]
  assign _T_2222 = _T_2218 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5091.6]
  assign V_121 = _T_2216 ? _T_2218 : _T_2222; // @[G128Multiplay.scala 46:7:@5084.4]
  assign _T_2224 = io_y[6]; // @[G128Multiplay.scala 37:16:@5095.4]
  assign _T_2227 = Z_121 ^ V_121; // @[G128Multiplay.scala 40:24:@5098.6]
  assign Z_122 = _T_2224 ? _T_2227 : Z_121; // @[G128Multiplay.scala 38:7:@5097.4]
  assign _T_2228 = V_121[0]; // @[G128Multiplay.scala 45:18:@5104.4]
  assign _T_2230 = _T_2228 == 1'h0; // @[G128Multiplay.scala 45:22:@5105.4]
  assign _T_2232 = V_121 >> 1'h1; // @[G128Multiplay.scala 48:24:@5107.6]
  assign _T_2236 = _T_2232 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5113.6]
  assign V_122 = _T_2230 ? _T_2232 : _T_2236; // @[G128Multiplay.scala 46:7:@5106.4]
  assign _T_2238 = io_y[5]; // @[G128Multiplay.scala 37:16:@5117.4]
  assign _T_2241 = Z_122 ^ V_122; // @[G128Multiplay.scala 40:24:@5120.6]
  assign Z_123 = _T_2238 ? _T_2241 : Z_122; // @[G128Multiplay.scala 38:7:@5119.4]
  assign _T_2242 = V_122[0]; // @[G128Multiplay.scala 45:18:@5126.4]
  assign _T_2244 = _T_2242 == 1'h0; // @[G128Multiplay.scala 45:22:@5127.4]
  assign _T_2246 = V_122 >> 1'h1; // @[G128Multiplay.scala 48:24:@5129.6]
  assign _T_2250 = _T_2246 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5135.6]
  assign V_123 = _T_2244 ? _T_2246 : _T_2250; // @[G128Multiplay.scala 46:7:@5128.4]
  assign _T_2252 = io_y[4]; // @[G128Multiplay.scala 37:16:@5139.4]
  assign _T_2255 = Z_123 ^ V_123; // @[G128Multiplay.scala 40:24:@5142.6]
  assign Z_124 = _T_2252 ? _T_2255 : Z_123; // @[G128Multiplay.scala 38:7:@5141.4]
  assign _T_2256 = V_123[0]; // @[G128Multiplay.scala 45:18:@5148.4]
  assign _T_2258 = _T_2256 == 1'h0; // @[G128Multiplay.scala 45:22:@5149.4]
  assign _T_2260 = V_123 >> 1'h1; // @[G128Multiplay.scala 48:24:@5151.6]
  assign _T_2264 = _T_2260 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5157.6]
  assign V_124 = _T_2258 ? _T_2260 : _T_2264; // @[G128Multiplay.scala 46:7:@5150.4]
  assign _T_2266 = io_y[3]; // @[G128Multiplay.scala 37:16:@5161.4]
  assign _T_2269 = Z_124 ^ V_124; // @[G128Multiplay.scala 40:24:@5164.6]
  assign Z_125 = _T_2266 ? _T_2269 : Z_124; // @[G128Multiplay.scala 38:7:@5163.4]
  assign _T_2270 = V_124[0]; // @[G128Multiplay.scala 45:18:@5170.4]
  assign _T_2272 = _T_2270 == 1'h0; // @[G128Multiplay.scala 45:22:@5171.4]
  assign _T_2274 = V_124 >> 1'h1; // @[G128Multiplay.scala 48:24:@5173.6]
  assign _T_2278 = _T_2274 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5179.6]
  assign V_125 = _T_2272 ? _T_2274 : _T_2278; // @[G128Multiplay.scala 46:7:@5172.4]
  assign _T_2280 = io_y[2]; // @[G128Multiplay.scala 37:16:@5183.4]
  assign _T_2283 = Z_125 ^ V_125; // @[G128Multiplay.scala 40:24:@5186.6]
  assign Z_126 = _T_2280 ? _T_2283 : Z_125; // @[G128Multiplay.scala 38:7:@5185.4]
  assign _T_2284 = V_125[0]; // @[G128Multiplay.scala 45:18:@5192.4]
  assign _T_2286 = _T_2284 == 1'h0; // @[G128Multiplay.scala 45:22:@5193.4]
  assign _T_2288 = V_125 >> 1'h1; // @[G128Multiplay.scala 48:24:@5195.6]
  assign _T_2292 = _T_2288 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5201.6]
  assign V_126 = _T_2286 ? _T_2288 : _T_2292; // @[G128Multiplay.scala 46:7:@5194.4]
  assign _T_2294 = io_y[1]; // @[G128Multiplay.scala 37:16:@5205.4]
  assign _T_2297 = Z_126 ^ V_126; // @[G128Multiplay.scala 40:24:@5208.6]
  assign Z_127 = _T_2294 ? _T_2297 : Z_126; // @[G128Multiplay.scala 38:7:@5207.4]
  assign _T_2298 = V_126[0]; // @[G128Multiplay.scala 45:18:@5214.4]
  assign _T_2300 = _T_2298 == 1'h0; // @[G128Multiplay.scala 45:22:@5215.4]
  assign _T_2302 = V_126 >> 1'h1; // @[G128Multiplay.scala 48:24:@5217.6]
  assign _T_2306 = _T_2302 ^ 128'he1000000000000000000000000000000; // @[G128Multiplay.scala 51:31:@5223.6]
  assign V_127 = _T_2300 ? _T_2302 : _T_2306; // @[G128Multiplay.scala 46:7:@5216.4]
  assign _T_2308 = io_y[0]; // @[G128Multiplay.scala 37:16:@5227.4]
  assign _T_2311 = Z_127 ^ V_127; // @[G128Multiplay.scala 40:24:@5230.6]
  assign Z_128 = _T_2308 ? _T_2311 : Z_127; // @[G128Multiplay.scala 38:7:@5229.4]
  assign io_out = Z_128;
endmodule
module pageswappergcm( // @[:@5251.2]
  input          clock, // @[:@5252.4]
  input          reset, // @[:@5253.4]
  input  [13:0]  io_mainMemio_addr, // @[:@5254.4]
  input          io_mainMemio_valid, // @[:@5254.4]
  input  [31:0]  io_mainMemio_wdata, // @[:@5254.4]
  input          io_mainMemio_we, // @[:@5254.4]
  input          io_mainMemio_en, // @[:@5254.4]
  output [31:0]  io_mainMemio_rdata, // @[:@5254.4]
  output         io_mainMemio_ready, // @[:@5254.4]
  output [13:0]  io_socMemio_addr, // @[:@5254.4]
  output [31:0]  io_socMemio_wdata, // @[:@5254.4]
  output         io_socMemio_we, // @[:@5254.4]
  output         io_socMemio_en, // @[:@5254.4]
  input  [31:0]  io_socMemio_rdata, // @[:@5254.4]
  input          io_socMemio_ready, // @[:@5254.4]
  output [10:0]  io_memio_addr, // @[:@5254.4]
  output [127:0] io_memio_wdata, // @[:@5254.4]
  output         io_memio_we, // @[:@5254.4]
  output         io_memio_en, // @[:@5254.4]
  input  [127:0] io_memio_rdata, // @[:@5254.4]
  input          io_memio_ready, // @[:@5254.4]
  output         io_err, // @[:@5254.4]
  output         io_currOutReady, // @[:@5254.4]
  output         io_finished // @[:@5254.4]
);
  wire  rndgenm_clock; // @[pageswappergcm.scala 28:23:@5256.4]
  wire  rndgenm_reset; // @[pageswappergcm.scala 28:23:@5256.4]
  wire [63:0] rndgenm_io_out; // @[pageswappergcm.scala 28:23:@5256.4]
  wire  rndgenm_io_en; // @[pageswappergcm.scala 28:23:@5256.4]
  wire  rndgenm_io_done; // @[pageswappergcm.scala 28:23:@5256.4]
  wire  cntrm_clock; // @[pageswappergcm.scala 29:23:@5259.4]
  wire  cntrm_io_get; // @[pageswappergcm.scala 29:23:@5259.4]
  wire [63:0] cntrm_io_out; // @[pageswappergcm.scala 29:23:@5259.4]
  wire  cntrm_io_reset; // @[pageswappergcm.scala 29:23:@5259.4]
  wire [63:0] cntrm_io_init; // @[pageswappergcm.scala 29:23:@5259.4]
  wire  vfm_clock; // @[pageswappergcm.scala 30:23:@5262.4]
  wire  vfm_reset; // @[pageswappergcm.scala 30:23:@5262.4]
  wire [127:0] vfm_io_rdata; // @[pageswappergcm.scala 30:23:@5262.4]
  wire [256:0] vfm_io_wdata; // @[pageswappergcm.scala 30:23:@5262.4]
  wire [4:0] vfm_io_addr; // @[pageswappergcm.scala 30:23:@5262.4]
  wire [2:0] vfm_io_cmd; // @[pageswappergcm.scala 30:23:@5262.4]
  wire  aesm_clock; // @[pageswappergcm.scala 31:23:@5265.4]
  wire  aesm_reset; // @[pageswappergcm.scala 31:23:@5265.4]
  wire [127:0] aesm_io_intVect; // @[pageswappergcm.scala 31:23:@5265.4]
  wire  aesm_io_newR; // @[pageswappergcm.scala 31:23:@5265.4]
  wire [127:0] aesm_io_out; // @[pageswappergcm.scala 31:23:@5265.4]
  wire [127:0] aesm_io_data; // @[pageswappergcm.scala 31:23:@5265.4]
  wire  aesm_io_en; // @[pageswappergcm.scala 31:23:@5265.4]
  wire [127:0] aesm_io_key; // @[pageswappergcm.scala 31:23:@5265.4]
  wire [127:0] gmultm_io_x; // @[pageswappergcm.scala 33:22:@5268.4]
  wire [127:0] gmultm_io_y; // @[pageswappergcm.scala 33:22:@5268.4]
  wire [127:0] gmultm_io_out; // @[pageswappergcm.scala 33:22:@5268.4]
  reg [127:0] h; // @[pageswappergcm.scala 34:18:@5271.4]
  reg [127:0] _RAND_0;
  reg [127:0] tag; // @[pageswappergcm.scala 35:20:@5272.4]
  reg [127:0] _RAND_1;
  reg [127:0] IVTag; // @[pageswappergcm.scala 36:22:@5273.4]
  reg [127:0] _RAND_2;
  reg [63:0] nonce; // @[pageswappergcm.scala 40:22:@5274.4]
  reg [63:0] _RAND_3;
  reg [127:0] curriv; // @[pageswappergcm.scala 41:23:@5275.4]
  reg [127:0] _RAND_4;
  reg [127:0] sessionIv; // @[pageswappergcm.scala 42:26:@5276.4]
  reg [127:0] _RAND_5;
  reg [127:0] sessionKey; // @[pageswappergcm.scala 44:27:@5277.4]
  reg [127:0] _RAND_6;
  reg [31:0] blockCounter; // @[pageswappergcm.scala 46:29:@5279.4]
  reg [31:0] _RAND_7;
  reg [127:0] currBlockBuff; // @[pageswappergcm.scala 47:30:@5280.4]
  reg [127:0] _RAND_8;
  reg [31:0] ConfReg_0; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_9;
  reg [31:0] ConfReg_1; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_10;
  reg [31:0] ConfReg_2; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_11;
  reg [31:0] ConfReg_3; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_12;
  reg [31:0] ConfReg_4; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_13;
  reg [31:0] ConfReg_5; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_14;
  reg [31:0] ConfReg_6; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_15;
  reg [31:0] ConfReg_7; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_16;
  reg [31:0] ConfReg_8; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_17;
  reg [31:0] ConfReg_9; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_18;
  reg [31:0] ConfReg_10; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_19;
  reg [31:0] ConfReg_11; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_20;
  reg [31:0] ConfReg_12; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_21;
  reg [31:0] ConfReg_13; // @[pageswappergcm.scala 96:20:@5312.4]
  reg [31:0] _RAND_22;
  reg [2:0] initState; // @[pageswappergcm.scala 108:26:@5327.4]
  reg [31:0] _RAND_23;
  reg [2:0] initStateNext; // @[pageswappergcm.scala 109:30:@5328.4]
  reg [31:0] _RAND_24;
  reg [2:0] poState; // @[pageswappergcm.scala 114:24:@5330.4]
  reg [31:0] _RAND_25;
  reg [1:0] cleanupState; // @[pageswappergcm.scala 118:29:@5333.4]
  reg [31:0] _RAND_26;
  reg [1:0] cleanupStateNext; // @[pageswappergcm.scala 119:33:@5334.4]
  reg [31:0] _RAND_27;
  reg [1:0] tagState; // @[pageswappergcm.scala 137:25:@5351.4]
  reg [31:0] _RAND_28;
  reg  tagUp; // @[pageswappergcm.scala 138:22:@5352.4]
  reg [31:0] _RAND_29;
  reg  encry; // @[pageswappergcm.scala 356:20:@5578.4]
  reg [31:0] _RAND_30;
  wire  start; // @[pageswappergcm.scala 125:25:@5337.4]
  wire [2:0] currOperation; // @[pageswappergcm.scala 126:33:@5338.4]
  wire  aesDone; // @[pageswappergcm.scala 128:27:@5339.4]
  wire [63:0] _T_216; // @[Cat.scala 30:58:@5340.4]
  wire [63:0] _T_217; // @[Cat.scala 30:58:@5341.4]
  wire [127:0] aesdecInput; // @[Cat.scala 30:58:@5342.4]
  wire  _T_219; // @[pageswappergcm.scala 130:37:@5343.4]
  wire  _T_221; // @[pageswappergcm.scala 130:63:@5344.4]
  wire  _T_222; // @[pageswappergcm.scala 130:46:@5345.4]
  wire [63:0] _T_223; // @[Cat.scala 30:58:@5346.4]
  wire [63:0] _T_224; // @[Cat.scala 30:58:@5347.4]
  wire [127:0] _T_225; // @[Cat.scala 30:58:@5348.4]
  wire [127:0] aesInOut; // @[pageswappergcm.scala 130:21:@5349.4]
  wire  moduleReady; // @[pageswappergcm.scala 134:31:@5350.4]
  wire [127:0] _T_238; // @[pageswappergcm.scala 145:82:@5358.4]
  wire [127:0] _T_239; // @[pageswappergcm.scala 145:102:@5359.4]
  wire [127:0] _T_240; // @[pageswappergcm.scala 145:24:@5360.4]
  wire [127:0] _T_241; // @[pageswappergcm.scala 144:20:@5361.4]
  wire [38:0] _GEN_425; // @[pageswappergcm.scala 147:31:@5362.4]
  wire [38:0] _T_242; // @[pageswappergcm.scala 147:31:@5362.4]
  wire [127:0] _GEN_426; // @[pageswappergcm.scala 147:37:@5363.4]
  wire [127:0] _T_243; // @[pageswappergcm.scala 147:37:@5363.4]
  wire  _T_244; // @[Mux.scala 46:19:@5364.4]
  wire [127:0] _T_245; // @[Mux.scala 46:16:@5365.4]
  wire  _T_246; // @[Mux.scala 46:19:@5366.4]
  wire [127:0] _T_247; // @[Mux.scala 46:16:@5367.4]
  wire  _T_248; // @[Mux.scala 46:19:@5368.4]
  wire [127:0] _T_249; // @[Mux.scala 46:16:@5369.4]
  wire  _T_251; // @[pageswappergcm.scala 151:28:@5371.4]
  wire  _T_253; // @[pageswappergcm.scala 151:53:@5372.4]
  wire [127:0] _T_255; // @[pageswappergcm.scala 151:64:@5373.4]
  wire [127:0] _T_256; // @[pageswappergcm.scala 151:43:@5374.4]
  wire [127:0] _T_257; // @[pageswappergcm.scala 151:15:@5375.4]
  wire  _T_260; // @[pageswappergcm.scala 155:27:@5378.4]
  wire [127:0] _T_261; // @[pageswappergcm.scala 155:18:@5379.4]
  wire  _T_263; // @[pageswappergcm.scala 156:33:@5380.4]
  wire [127:0] _T_264; // @[pageswappergcm.scala 156:71:@5381.4]
  wire [127:0] _T_265; // @[pageswappergcm.scala 156:19:@5382.4]
  wire [127:0] _T_267; // @[Mux.scala 46:16:@5384.4]
  wire [127:0] _T_269; // @[Mux.scala 46:16:@5386.4]
  wire  _T_270; // @[pageswappergcm.scala 160:31:@5388.4]
  wire  _T_274; // @[pageswappergcm.scala 173:56:@5392.4]
  wire  _T_275; // @[pageswappergcm.scala 173:43:@5393.4]
  wire  _T_279; // @[pageswappergcm.scala 175:48:@5398.4]
  wire [63:0] _T_281; // @[pageswappergcm.scala 175:23:@5399.4]
  wire  cond1; // @[pageswappergcm.scala 177:24:@5401.4]
  wire  cond2; // @[pageswappergcm.scala 178:28:@5402.4]
  wire  _T_283; // @[pageswappergcm.scala 180:35:@5404.4]
  wire  _T_284; // @[pageswappergcm.scala 180:48:@5405.4]
  wire  _T_285; // @[pageswappergcm.scala 180:22:@5406.4]
  wire  cond4; // @[pageswappergcm.scala 180:60:@5407.4]
  wire  _T_287; // @[pageswappergcm.scala 181:48:@5409.4]
  wire  _T_288; // @[pageswappergcm.scala 181:66:@5410.4]
  wire  _T_289; // @[pageswappergcm.scala 181:22:@5411.4]
  wire  cond5; // @[pageswappergcm.scala 181:78:@5412.4]
  wire  _T_290; // @[pageswappergcm.scala 183:26:@5413.4]
  wire  _T_291; // @[pageswappergcm.scala 183:53:@5414.4]
  wire  _T_292; // @[pageswappergcm.scala 183:37:@5415.4]
  wire  newc24; // @[pageswappergcm.scala 183:64:@5416.4]
  wire  _T_298; // @[Mux.scala 46:19:@5417.4]
  wire  _T_299; // @[Mux.scala 46:16:@5418.4]
  wire  _T_300; // @[Mux.scala 46:19:@5419.4]
  wire  _T_301; // @[Mux.scala 46:16:@5420.4]
  wire  _T_302; // @[Mux.scala 46:19:@5421.4]
  wire  _T_303; // @[Mux.scala 46:16:@5422.4]
  wire  _T_304; // @[Mux.scala 46:19:@5423.4]
  wire  cond; // @[Mux.scala 46:16:@5424.4]
  wire  newC; // @[pageswappergcm.scala 192:14:@5426.4]
  wire  _T_311; // @[pageswappergcm.scala 206:44:@5428.4]
  wire [1:0] _T_314; // @[pageswappergcm.scala 206:30:@5429.4]
  wire  _T_316; // @[Mux.scala 46:19:@5430.4]
  wire [2:0] _T_317; // @[Mux.scala 46:16:@5431.4]
  wire  _T_318; // @[Mux.scala 46:19:@5432.4]
  wire [2:0] x1; // @[Mux.scala 46:16:@5433.4]
  wire  _T_325; // @[Mux.scala 46:19:@5434.4]
  wire [1:0] _T_326; // @[Mux.scala 46:16:@5435.4]
  wire  _T_327; // @[Mux.scala 46:19:@5436.4]
  wire [2:0] _T_328; // @[Mux.scala 46:16:@5437.4]
  wire  _T_330; // @[Mux.scala 46:19:@5438.4]
  wire [2:0] x3; // @[Mux.scala 46:16:@5441.4]
  wire [1:0] _T_341; // @[Mux.scala 46:16:@5445.4]
  wire  _T_342; // @[Mux.scala 46:19:@5446.4]
  wire [1:0] x2; // @[Mux.scala 46:16:@5447.4]
  wire  _T_350; // @[pageswappergcm.scala 231:47:@5450.4]
  wire [1:0] _T_353; // @[pageswappergcm.scala 231:32:@5451.4]
  wire  _T_355; // @[pageswappergcm.scala 232:43:@5452.4]
  wire [1:0] _T_358; // @[pageswappergcm.scala 232:29:@5453.4]
  wire  _T_359; // @[Mux.scala 46:19:@5454.4]
  wire [1:0] _T_360; // @[Mux.scala 46:16:@5455.4]
  wire  _T_361; // @[Mux.scala 46:19:@5456.4]
  wire [1:0] _T_362; // @[Mux.scala 46:16:@5457.4]
  wire [1:0] x4; // @[Mux.scala 46:16:@5459.4]
  wire [1:0] _T_370; // @[Mux.scala 46:16:@5461.4]
  wire [2:0] _T_372; // @[Mux.scala 46:16:@5463.4]
  wire [2:0] _T_374; // @[Mux.scala 46:16:@5465.4]
  wire [2:0] _T_376; // @[Mux.scala 46:16:@5467.4]
  wire  _T_378; // @[pageswappergcm.scala 250:27:@5469.4]
  wire [31:0] _T_380; // @[pageswappergcm.scala 250:18:@5470.4]
  wire [32:0] _T_386; // @[pageswappergcm.scala 254:70:@5472.4]
  wire [32:0] _T_387; // @[pageswappergcm.scala 254:70:@5473.4]
  wire [31:0] _T_388; // @[pageswappergcm.scala 254:70:@5474.4]
  wire [31:0] _T_389; // @[pageswappergcm.scala 254:35:@5475.4]
  wire [31:0] _T_391; // @[Mux.scala 46:16:@5477.4]
  wire [31:0] _T_393; // @[Mux.scala 46:16:@5479.4]
  wire [31:0] _T_395; // @[Mux.scala 46:16:@5481.4]
  wire [382:0] _GEN_427; // @[pageswappergcm.scala 264:40:@5483.4]
  wire [382:0] _T_400; // @[pageswappergcm.scala 264:40:@5483.4]
  wire [382:0] _GEN_428; // @[pageswappergcm.scala 264:49:@5484.4]
  wire [382:0] _T_401; // @[pageswappergcm.scala 264:49:@5484.4]
  wire [383:0] _T_402; // @[Cat.scala 30:58:@5485.4]
  wire [383:0] _T_408; // @[Cat.scala 30:58:@5488.4]
  wire [382:0] _GEN_433; // @[pageswappergcm.scala 267:39:@5492.4]
  wire [382:0] _T_418; // @[pageswappergcm.scala 267:39:@5492.4]
  wire [382:0] _T_419; // @[pageswappergcm.scala 267:48:@5493.4]
  wire [383:0] _T_420; // @[Cat.scala 30:58:@5494.4]
  wire [383:0] _T_422; // @[Mux.scala 46:16:@5496.4]
  wire [383:0] _T_424; // @[Mux.scala 46:16:@5498.4]
  wire [383:0] _T_426; // @[Mux.scala 46:16:@5500.4]
  wire [383:0] _T_428; // @[Mux.scala 46:16:@5502.4]
  wire [190:0] _GEN_435; // @[pageswappergcm.scala 277:30:@5504.4]
  wire [190:0] _T_430; // @[pageswappergcm.scala 277:30:@5504.4]
  wire [190:0] _GEN_436; // @[pageswappergcm.scala 277:38:@5505.4]
  wire [190:0] _T_431; // @[pageswappergcm.scala 277:38:@5505.4]
  wire [190:0] cv13; // @[pageswappergcm.scala 277:17:@5506.4]
  wire  _T_435; // @[pageswappergcm.scala 278:37:@5509.4]
  wire  _T_436; // @[pageswappergcm.scala 279:18:@5510.4]
  wire [128:0] _T_438; // @[pageswappergcm.scala 279:40:@5511.4]
  wire [127:0] _T_439; // @[pageswappergcm.scala 279:40:@5512.4]
  wire [127:0] _T_440; // @[pageswappergcm.scala 279:8:@5513.4]
  wire [127:0] cv2; // @[pageswappergcm.scala 278:17:@5514.4]
  wire [127:0] _T_446; // @[Mux.scala 46:16:@5516.4]
  wire [127:0] _T_448; // @[Mux.scala 46:16:@5518.4]
  wire [190:0] _T_450; // @[Mux.scala 46:16:@5520.4]
  wire [190:0] xcv; // @[Mux.scala 46:16:@5522.4]
  wire [190:0] _T_454; // @[pageswappergcm.scala 298:20:@5525.4]
  wire [127:0] _T_460; // @[pageswappergcm.scala 300:20:@5529.4]
  wire  _T_462; // @[pageswappergcm.scala 301:30:@5530.4]
  wire  _T_465; // @[pageswappergcm.scala 301:41:@5532.4]
  wire [127:0] _T_466; // @[pageswappergcm.scala 301:20:@5533.4]
  wire [127:0] _T_468; // @[Mux.scala 46:16:@5535.4]
  wire [127:0] _T_470; // @[Mux.scala 46:16:@5537.4]
  wire [190:0] _T_472; // @[Mux.scala 46:16:@5539.4]
  wire [190:0] _T_474; // @[Mux.scala 46:16:@5541.4]
  wire  _T_476; // @[pageswappergcm.scala 313:31:@5543.4]
  wire  bcg1; // @[pageswappergcm.scala 313:17:@5545.4]
  wire  _T_480; // @[pageswappergcm.scala 314:31:@5546.4]
  wire  bcg2; // @[pageswappergcm.scala 314:17:@5548.4]
  wire  _T_489; // @[Mux.scala 46:16:@5550.4]
  wire  _T_491; // @[Mux.scala 46:16:@5552.4]
  wire  _T_493; // @[Mux.scala 46:16:@5554.4]
  wire  _T_495; // @[Mux.scala 46:16:@5556.4]
  wire  _T_497; // @[pageswappergcm.scala 340:24:@5558.4]
  wire  _T_498; // @[pageswappergcm.scala 341:28:@5560.4]
  wire [127:0] _T_503; // @[pageswappergcm.scala 346:43:@5564.4]
  wire [127:0] _T_504; // @[pageswappergcm.scala 346:18:@5565.4]
  wire [127:0] _T_508; // @[pageswappergcm.scala 347:18:@5567.4]
  wire [127:0] _T_512; // @[Mux.scala 46:16:@5569.4]
  wire [127:0] _T_514; // @[Mux.scala 46:16:@5571.4]
  wire [127:0] _T_516; // @[Mux.scala 46:16:@5573.4]
  wire [127:0] cb; // @[Mux.scala 46:16:@5575.4]
  wire  _T_522; // @[pageswappergcm.scala 357:46:@5580.4]
  wire  _T_524; // @[pageswappergcm.scala 357:14:@5582.4]
  wire [127:0] _T_528; // @[pageswappergcm.scala 359:25:@5586.4]
  wire [127:0] _T_533; // @[pageswappergcm.scala 363:29:@5589.4]
  wire [127:0] _T_543; // @[pageswappergcm.scala 365:29:@5593.4]
  wire [127:0] _T_550; // @[Mux.scala 46:16:@5597.4]
  wire [127:0] _T_552; // @[Mux.scala 46:16:@5599.4]
  wire [127:0] _T_554; // @[Mux.scala 46:16:@5601.4]
  wire [127:0] _T_556; // @[Mux.scala 46:16:@5603.4]
  wire  socmselect; // @[pageswappergcm.scala 387:38:@5622.4]
  wire  _T_583; // @[pageswappergcm.scala 388:44:@5623.4]
  wire [14:0] _T_586; // @[pageswappergcm.scala 388:123:@5624.4]
  wire [13:0] _T_587; // @[pageswappergcm.scala 388:123:@5625.4]
  wire  _T_588; // @[pageswappergcm.scala 388:94:@5626.4]
  wire  validConfAddress; // @[pageswappergcm.scala 388:73:@5627.4]
  wire  _T_590; // @[pageswappergcm.scala 393:45:@5630.4]
  wire  _T_591; // @[pageswappergcm.scala 393:54:@5631.4]
  wire  _T_598; // @[pageswappergcm.scala 394:29:@5636.4]
  wire  _T_603; // @[pageswappergcm.scala 395:29:@5640.4]
  wire [3:0] confaddr; // @[pageswappergcm.scala 398:35:@5642.4]
  wire [31:0] _T_811; // @[pageswappergcm.scala 635:42:@5848.20]
  wire [31:0] _GEN_121; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_158; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_175; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_191; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_206; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_330; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_351; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] ConfRegWire_1; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _T_810; // @[pageswappergcm.scala 634:42:@5846.20]
  wire [31:0] _GEN_120; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_157; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_174; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_190; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_205; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_329; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_350; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] ConfRegWire_0; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_4; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _T_812; // @[pageswappergcm.scala 636:42:@5850.20]
  wire [31:0] _GEN_122; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_159; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_176; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_192; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_207; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_331; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_352; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] ConfRegWire_2; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_5; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _T_813; // @[pageswappergcm.scala 637:42:@5852.20]
  wire [31:0] _GEN_123; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_160; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_177; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_193; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_208; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_332; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_353; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] ConfRegWire_3; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_6; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_7; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_8; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_9; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_10; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_11; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_12; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_13; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_14; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_15; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _GEN_16; // @[pageswappergcm.scala 412:29:@5645.4]
  wire [31:0] _T_608; // @[pageswappergcm.scala 412:29:@5645.4]
  wire  _T_611; // @[pageswappergcm.scala 416:55:@5647.4]
  wire  _T_616; // @[pageswappergcm.scala 417:41:@5649.4]
  wire  _T_618; // @[Mux.scala 46:16:@5651.4]
  wire  _T_619; // @[Mux.scala 46:19:@5652.4]
  wire  _T_620; // @[Mux.scala 46:16:@5653.4]
  wire  _T_625; // @[Mux.scala 46:19:@5656.4]
  wire [31:0] confMask; // @[Mux.scala 46:16:@5657.4]
  wire  _T_627; // @[pageswappergcm.scala 437:42:@5658.4]
  wire  _T_629; // @[pageswappergcm.scala 437:69:@5659.4]
  wire  _T_630; // @[pageswappergcm.scala 437:51:@5660.4]
  wire  _T_631; // @[pageswappergcm.scala 437:90:@5661.4]
  wire  pindataReady; // @[pageswappergcm.scala 437:25:@5662.4]
  wire  _T_638; // @[pageswappergcm.scala 438:91:@5666.4]
  wire  poutdataReady; // @[pageswappergcm.scala 438:26:@5667.4]
  wire  _T_641; // @[pageswappergcm.scala 447:14:@5671.6]
  wire  _T_642; // @[pageswappergcm.scala 447:26:@5672.6]
  wire [31:0] _T_643; // @[pageswappergcm.scala 451:48:@5675.10]
  wire [31:0] _T_644; // @[pageswappergcm.scala 451:45:@5676.10]
  wire  _T_646; // @[pageswappergcm.scala 455:35:@5677.10]
  wire  _T_647; // @[pageswappergcm.scala 456:19:@5678.10]
  wire [31:0] _GEN_17; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_18; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_19; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_20; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_21; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_22; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_23; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_24; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_25; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_26; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_27; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_28; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_29; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _T_656; // @[pageswappergcm.scala 463:85:@5682.12]
  wire [31:0] _GEN_30; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_31; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_32; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_35; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_36; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_37; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_38; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_39; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_40; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_41; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_42; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_43; // @[pageswappergcm.scala 463:50:@5683.12]
  wire [31:0] _GEN_44; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_45; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_46; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_49; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_50; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_51; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_52; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_53; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_54; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_55; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_56; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_57; // @[pageswappergcm.scala 472:50:@5687.12]
  wire [31:0] _GEN_58; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_59; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_60; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_63; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_64; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_65; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_66; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_67; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_68; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_69; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_70; // @[pageswappergcm.scala 457:14:@5679.10]
  wire [31:0] _GEN_71; // @[pageswappergcm.scala 457:14:@5679.10]
  wire  _T_667; // @[pageswappergcm.scala 476:95:@5692.10]
  wire  _T_668; // @[pageswappergcm.scala 476:77:@5693.10]
  wire  _T_671; // @[pageswappergcm.scala 476:132:@5695.10]
  wire  _T_672; // @[pageswappergcm.scala 476:105:@5696.10]
  wire [7:0] _T_675; // @[pageswappergcm.scala 479:47:@5698.12]
  wire [31:0] _GEN_437; // @[pageswappergcm.scala 479:41:@5699.12]
  wire [31:0] _T_676; // @[pageswappergcm.scala 479:41:@5699.12]
  wire [31:0] _GEN_72; // @[pageswappergcm.scala 478:14:@5697.10]
  wire [31:0] _GEN_73; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_74; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_75; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_78; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_79; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_80; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_81; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_82; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_83; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_84; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_85; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_86; // @[pageswappergcm.scala 450:12:@5674.8]
  wire [31:0] _GEN_87; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_88; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_89; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_92; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_93; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_94; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_95; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_96; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_97; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_98; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_99; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_100; // @[pageswappergcm.scala 448:9:@5673.6]
  wire [31:0] _GEN_101; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_102; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_103; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_106; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_107; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_108; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_109; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_110; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_111; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_112; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_113; // @[pageswappergcm.scala 445:3:@5670.4]
  wire [31:0] _GEN_114; // @[pageswappergcm.scala 445:3:@5670.4]
  wire  vfNotFull; // @[pageswappergcm.scala 498:34:@5707.4]
  wire  _T_681; // @[pageswappergcm.scala 502:42:@5709.4]
  wire [127:0] _T_683; // @[pageswappergcm.scala 502:22:@5710.4]
  wire [31:0] _T_686; // @[Mux.scala 46:16:@5712.4]
  wire [127:0] conf3; // @[Mux.scala 46:16:@5714.4]
  wire [127:0] _T_689; // @[pageswappergcm.scala 505:22:@5716.4]
  wire  _T_693; // @[pageswappergcm.scala 511:44:@5719.4]
  wire  _T_694; // @[pageswappergcm.scala 511:41:@5720.4]
  wire [31:0] _T_696; // @[pageswappergcm.scala 511:68:@5721.4]
  wire [31:0] _T_697; // @[pageswappergcm.scala 511:20:@5722.4]
  wire [31:0] conf4; // @[Mux.scala 46:16:@5724.4]
  wire [31:0] _T_700; // @[pageswappergcm.scala 513:22:@5726.4]
  wire  _T_713; // @[Mux.scala 46:16:@5733.4]
  wire  mmenvalid; // @[Mux.scala 46:16:@5735.4]
  wire [10:0] _T_720; // @[pageswappergcm.scala 533:27:@5741.4]
  wire [31:0] _GEN_438; // @[pageswappergcm.scala 533:63:@5745.4]
  wire [32:0] _T_725; // @[pageswappergcm.scala 533:63:@5745.4]
  wire [31:0] addr2; // @[pageswappergcm.scala 533:63:@5746.4]
  wire [32:0] _T_727; // @[pageswappergcm.scala 536:63:@5748.4]
  wire [31:0] addr1; // @[pageswappergcm.scala 536:63:@5749.4]
  wire [31:0] _T_732; // @[pageswappergcm.scala 541:19:@5751.4]
  wire [31:0] _T_736; // @[pageswappergcm.scala 542:19:@5753.4]
  wire [31:0] _T_738; // @[Mux.scala 46:16:@5755.4]
  wire [31:0] addr; // @[Mux.scala 46:16:@5757.4]
  wire  _T_743; // @[pageswappergcm.scala 546:48:@5761.4]
  wire [127:0] _T_748; // @[pageswappergcm.scala 546:25:@5765.4]
  wire [2:0] nPoState; // @[pageswappergcm.scala 552:21:@5769.4]
  wire [2:0] _T_751; // @[pageswappergcm.scala 559:40:@5770.4]
  wire [2:0] _T_752; // @[pageswappergcm.scala 559:23:@5771.4]
  wire [2:0] _T_753; // @[pageswappergcm.scala 560:47:@5772.4]
  wire [2:0] _T_754; // @[pageswappergcm.scala 560:29:@5773.4]
  wire [2:0] _T_757; // @[pageswappergcm.scala 561:50:@5775.4]
  wire [2:0] _T_758; // @[pageswappergcm.scala 561:24:@5776.4]
  wire [2:0] _T_761; // @[pageswappergcm.scala 562:24:@5778.4]
  wire [2:0] _T_763; // @[Mux.scala 46:16:@5780.4]
  wire [2:0] _T_765; // @[Mux.scala 46:16:@5782.4]
  wire  _T_766; // @[Mux.scala 46:19:@5783.4]
  wire [2:0] _T_767; // @[Mux.scala 46:16:@5784.4]
  wire [2:0] _T_769; // @[Mux.scala 46:16:@5786.4]
  wire [2:0] _T_771; // @[Mux.scala 46:16:@5788.4]
  wire [2:0] pos13; // @[Mux.scala 46:16:@5790.4]
  wire  _T_773; // @[pageswappergcm.scala 566:28:@5791.4]
  wire [2:0] _T_774; // @[pageswappergcm.scala 566:21:@5792.4]
  wire [34:0] _T_785; // @[pageswappergcm.scala 588:49:@5804.12]
  wire [34:0] _T_786; // @[pageswappergcm.scala 588:38:@5805.12]
  wire [34:0] _GEN_440; // @[pageswappergcm.scala 588:36:@5806.12]
  wire [34:0] _T_787; // @[pageswappergcm.scala 588:36:@5806.12]
  wire [31:0] _GEN_115; // @[pageswappergcm.scala 595:13:@5813.14]
  wire [1:0] _GEN_116; // @[pageswappergcm.scala 595:13:@5813.14]
  wire [3:0] _T_796; // @[pageswappergcm.scala 604:46:@5821.16]
  wire [3:0] _T_797; // @[pageswappergcm.scala 604:41:@5822.16]
  wire [31:0] _GEN_441; // @[pageswappergcm.scala 604:38:@5823.16]
  wire [31:0] _T_798; // @[pageswappergcm.scala 604:38:@5823.16]
  wire [32:0] _T_802; // @[pageswappergcm.scala 616:46:@5828.20]
  wire [31:0] _T_803; // @[pageswappergcm.scala 616:46:@5829.20]
  wire [31:0] _GEN_117; // @[pageswappergcm.scala 614:15:@5827.18]
  wire [31:0] _GEN_118; // @[pageswappergcm.scala 621:13:@5835.18]
  wire [31:0] _GEN_119; // @[pageswappergcm.scala 606:13:@5826.16]
  wire [31:0] _GEN_442; // @[pageswappergcm.scala 655:38:@5864.20]
  wire [31:0] _T_822; // @[pageswappergcm.scala 655:38:@5864.20]
  wire [31:0] _GEN_124; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_125; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_126; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_127; // @[pageswappergcm.scala 632:11:@5845.18]
  wire  _GEN_128; // @[pageswappergcm.scala 632:11:@5845.18]
  wire [31:0] _GEN_129; // @[pageswappergcm.scala 632:11:@5845.18]
  wire  _T_823; // @[pageswappergcm.scala 683:28:@5869.18]
  wire [38:0] _T_827; // @[pageswappergcm.scala 691:55:@5873.22]
  wire [38:0] _T_828; // @[pageswappergcm.scala 691:44:@5874.22]
  wire [38:0] _GEN_443; // @[pageswappergcm.scala 691:42:@5875.22]
  wire [38:0] _T_829; // @[pageswappergcm.scala 691:42:@5875.22]
  wire [38:0] _GEN_130; // @[pageswappergcm.scala 689:15:@5872.20]
  wire  _T_835; // @[pageswappergcm.scala 708:37:@5888.24]
  wire [31:0] _T_840; // @[pageswappergcm.scala 715:41:@5896.28]
  wire [38:0] _T_843; // @[pageswappergcm.scala 716:53:@5898.28]
  wire [38:0] _T_844; // @[pageswappergcm.scala 716:41:@5899.28]
  wire [31:0] _GEN_131; // @[pageswappergcm.scala 713:12:@5895.26]
  wire [38:0] _GEN_132; // @[pageswappergcm.scala 713:12:@5895.26]
  wire [1:0] _GEN_133; // @[pageswappergcm.scala 713:12:@5895.26]
  wire [31:0] _GEN_134; // @[pageswappergcm.scala 713:12:@5895.26]
  wire [1:0] _GEN_135; // @[pageswappergcm.scala 713:12:@5895.26]
  wire [1:0] _GEN_136; // @[pageswappergcm.scala 709:12:@5889.24]
  wire [1:0] _GEN_137; // @[pageswappergcm.scala 709:12:@5889.24]
  wire [31:0] _GEN_138; // @[pageswappergcm.scala 709:12:@5889.24]
  wire [38:0] _GEN_139; // @[pageswappergcm.scala 709:12:@5889.24]
  wire [31:0] _GEN_140; // @[pageswappergcm.scala 709:12:@5889.24]
  wire [1:0] _GEN_141; // @[pageswappergcm.scala 704:12:@5884.22]
  wire [1:0] _GEN_142; // @[pageswappergcm.scala 704:12:@5884.22]
  wire [31:0] _GEN_143; // @[pageswappergcm.scala 704:12:@5884.22]
  wire [38:0] _GEN_144; // @[pageswappergcm.scala 704:12:@5884.22]
  wire [31:0] _GEN_145; // @[pageswappergcm.scala 704:12:@5884.22]
  wire [1:0] _GEN_146; // @[pageswappergcm.scala 697:9:@5881.20]
  wire [1:0] _GEN_147; // @[pageswappergcm.scala 697:9:@5881.20]
  wire [31:0] _GEN_148; // @[pageswappergcm.scala 697:9:@5881.20]
  wire [38:0] _GEN_149; // @[pageswappergcm.scala 697:9:@5881.20]
  wire [31:0] _GEN_150; // @[pageswappergcm.scala 697:9:@5881.20]
  wire  _GEN_151; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [38:0] _GEN_152; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [1:0] _GEN_153; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [1:0] _GEN_154; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [31:0] _GEN_155; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [31:0] _GEN_156; // @[pageswappergcm.scala 684:9:@5870.18]
  wire [31:0] _GEN_161; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_162; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_163; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_164; // @[pageswappergcm.scala 629:9:@5844.16]
  wire  _GEN_165; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [38:0] _GEN_166; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [1:0] _GEN_167; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [1:0] _GEN_168; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_169; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [31:0] _GEN_170; // @[pageswappergcm.scala 629:9:@5844.16]
  wire [38:0] _GEN_171; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_172; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [1:0] _GEN_173; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_178; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_179; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_180; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_181; // @[pageswappergcm.scala 602:9:@5820.14]
  wire  _GEN_182; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [1:0] _GEN_183; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_184; // @[pageswappergcm.scala 602:9:@5820.14]
  wire [31:0] _GEN_185; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [1:0] _GEN_186; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [38:0] _GEN_187; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_188; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [1:0] _GEN_189; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_194; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_195; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_196; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_197; // @[pageswappergcm.scala 591:9:@5811.12]
  wire  _GEN_198; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [31:0] _GEN_199; // @[pageswappergcm.scala 591:9:@5811.12]
  wire [38:0] _GEN_200; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_201; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [1:0] _GEN_202; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_203; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [1:0] _GEN_204; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_209; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_210; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_211; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_212; // @[pageswappergcm.scala 586:9:@5803.10]
  wire  _GEN_213; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_214; // @[pageswappergcm.scala 586:9:@5803.10]
  wire [31:0] _GEN_215; // @[pageswappergcm.scala 736:13:@5924.14]
  wire [1:0] _GEN_216; // @[pageswappergcm.scala 736:13:@5924.14]
  wire [38:0] _T_868; // @[pageswappergcm.scala 749:53:@5938.20]
  wire [38:0] _T_869; // @[pageswappergcm.scala 749:42:@5939.20]
  wire [38:0] _T_870; // @[pageswappergcm.scala 749:40:@5940.20]
  wire [38:0] _GEN_217; // @[pageswappergcm.scala 748:13:@5937.18]
  wire [2:0] _GEN_218; // @[pageswappergcm.scala 748:13:@5937.18]
  wire [31:0] _GEN_219; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [31:0] _GEN_220; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [31:0] _GEN_221; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [31:0] _GEN_222; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [2:0] _GEN_223; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [31:0] _GEN_225; // @[pageswappergcm.scala 755:13:@5948.20]
  wire [32:0] _T_890; // @[pageswappergcm.scala 776:33:@5973.22]
  wire [32:0] _T_891; // @[pageswappergcm.scala 776:33:@5974.22]
  wire [31:0] _T_892; // @[pageswappergcm.scala 776:33:@5975.22]
  wire  _T_894; // @[pageswappergcm.scala 776:39:@5976.22]
  wire  _T_901; // @[pageswappergcm.scala 792:45:@5987.28]
  wire [2:0] _GEN_226; // @[pageswappergcm.scala 793:21:@5988.28]
  wire [2:0] _GEN_227; // @[pageswappergcm.scala 790:19:@5983.26]
  wire [2:0] _GEN_229; // @[pageswappergcm.scala 782:17:@5982.24]
  wire [2:0] _GEN_230; // @[pageswappergcm.scala 777:15:@5977.22]
  wire [38:0] _T_926; // @[pageswappergcm.scala 829:59:@6034.30]
  wire  _T_929; // @[pageswappergcm.scala 842:30:@6040.30]
  wire [31:0] _T_932; // @[pageswappergcm.scala 844:42:@6043.32]
  wire [31:0] _T_934; // @[pageswappergcm.scala 847:42:@6047.32]
  wire [31:0] _GEN_231; // @[pageswappergcm.scala 843:15:@6041.30]
  wire [38:0] _GEN_233; // @[pageswappergcm.scala 826:12:@6027.28]
  wire [2:0] _GEN_234; // @[pageswappergcm.scala 826:12:@6027.28]
  wire [31:0] _GEN_238; // @[pageswappergcm.scala 826:12:@6027.28]
  wire [38:0] _GEN_242; // @[pageswappergcm.scala 822:12:@6021.26]
  wire [2:0] _GEN_243; // @[pageswappergcm.scala 822:12:@6021.26]
  wire [31:0] _GEN_245; // @[pageswappergcm.scala 822:12:@6021.26]
  wire [38:0] _GEN_249; // @[pageswappergcm.scala 817:12:@6016.24]
  wire [2:0] _GEN_250; // @[pageswappergcm.scala 817:12:@6016.24]
  wire [31:0] _GEN_252; // @[pageswappergcm.scala 817:12:@6016.24]
  wire [38:0] _GEN_256; // @[pageswappergcm.scala 810:11:@6013.22]
  wire [2:0] _GEN_257; // @[pageswappergcm.scala 810:11:@6013.22]
  wire [31:0] _GEN_259; // @[pageswappergcm.scala 810:11:@6013.22]
  wire [38:0] _GEN_260; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [2:0] _GEN_261; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [1:0] _GEN_262; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [1:0] _GEN_263; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [31:0] _GEN_264; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [31:0] _GEN_265; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [31:0] _GEN_266; // @[pageswappergcm.scala 774:11:@5968.20]
  wire [31:0] _GEN_267; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_268; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_269; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_270; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [2:0] _GEN_271; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [38:0] _GEN_272; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_273; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [1:0] _GEN_274; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [1:0] _GEN_275; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_276; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [31:0] _GEN_277; // @[pageswappergcm.scala 753:11:@5947.18]
  wire [38:0] _GEN_278; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [2:0] _GEN_279; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_280; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_281; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_282; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_283; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_284; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [1:0] _GEN_285; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [1:0] _GEN_286; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_287; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [31:0] _GEN_288; // @[pageswappergcm.scala 746:11:@5936.16]
  wire [2:0] _GEN_289; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [38:0] _GEN_290; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_291; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_292; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_293; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_294; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_295; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [1:0] _GEN_296; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [1:0] _GEN_297; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_298; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [31:0] _GEN_299; // @[pageswappergcm.scala 743:11:@5931.14]
  wire [2:0] _GEN_300; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [38:0] _GEN_301; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_302; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [1:0] _GEN_303; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_304; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_305; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_306; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_307; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_308; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [1:0] _GEN_309; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_310; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [31:0] _GEN_311; // @[pageswappergcm.scala 731:11:@5917.12]
  wire [2:0] _GEN_312; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [38:0] _GEN_313; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_314; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [1:0] _GEN_315; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_316; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_317; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_318; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_319; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_320; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [1:0] _GEN_321; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_322; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [31:0] _GEN_323; // @[pageswappergcm.scala 729:7:@5915.10]
  wire [38:0] _GEN_324; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_325; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [1:0] _GEN_326; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_327; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [1:0] _GEN_328; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_333; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_334; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_335; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_336; // @[pageswappergcm.scala 583:7:@5801.8]
  wire  _GEN_337; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_338; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [2:0] _GEN_339; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_340; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_341; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_342; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_343; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [31:0] _GEN_344; // @[pageswappergcm.scala 583:7:@5801.8]
  wire [38:0] _GEN_345; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_346; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [1:0] _GEN_347; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_348; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [1:0] _GEN_349; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_354; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_355; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_356; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_357; // @[pageswappergcm.scala 580:5:@5797.6]
  wire  _GEN_358; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_359; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [2:0] _GEN_360; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_361; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_362; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_363; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_364; // @[pageswappergcm.scala 580:5:@5797.6]
  wire [31:0] _GEN_365; // @[pageswappergcm.scala 580:5:@5797.6]
  wire  _T_937; // @[pageswappergcm.scala 862:20:@6060.6]
  wire  _T_938; // @[pageswappergcm.scala 865:26:@6065.8]
  wire [63:0] _GEN_366; // @[pageswappergcm.scala 868:11:@6067.10]
  wire [2:0] _GEN_367; // @[pageswappergcm.scala 868:11:@6067.10]
  wire  _T_939; // @[pageswappergcm.scala 872:26:@6073.10]
  wire [127:0] _GEN_368; // @[pageswappergcm.scala 875:11:@6075.12]
  wire [2:0] _GEN_369; // @[pageswappergcm.scala 875:11:@6075.12]
  wire  _T_940; // @[pageswappergcm.scala 879:26:@6081.12]
  wire [190:0] _GEN_450; // @[pageswappergcm.scala 883:51:@6084.16]
  wire [190:0] _T_942; // @[pageswappergcm.scala 883:51:@6084.16]
  wire [190:0] _GEN_451; // @[pageswappergcm.scala 883:34:@6085.16]
  wire [190:0] _T_943; // @[pageswappergcm.scala 883:34:@6085.16]
  wire [190:0] _GEN_370; // @[pageswappergcm.scala 882:11:@6083.14]
  wire [2:0] _GEN_371; // @[pageswappergcm.scala 882:11:@6083.14]
  wire [2:0] _GEN_372; // @[pageswappergcm.scala 890:9:@6093.16]
  wire [1:0] _T_948; // @[pageswappergcm.scala 903:46:@6102.20]
  wire [31:0] _GEN_452; // @[pageswappergcm.scala 903:40:@6103.20]
  wire [31:0] _T_949; // @[pageswappergcm.scala 903:40:@6103.20]
  wire [127:0] _GEN_373; // @[pageswappergcm.scala 896:11:@6100.18]
  wire [31:0] _GEN_374; // @[pageswappergcm.scala 896:11:@6100.18]
  wire [2:0] _GEN_375; // @[pageswappergcm.scala 896:11:@6100.18]
  wire [127:0] _GEN_376; // @[pageswappergcm.scala 894:6:@6099.16]
  wire [31:0] _GEN_377; // @[pageswappergcm.scala 894:6:@6099.16]
  wire [2:0] _GEN_378; // @[pageswappergcm.scala 894:6:@6099.16]
  wire [2:0] _GEN_379; // @[pageswappergcm.scala 888:6:@6092.14]
  wire [127:0] _GEN_380; // @[pageswappergcm.scala 888:6:@6092.14]
  wire [31:0] _GEN_381; // @[pageswappergcm.scala 888:6:@6092.14]
  wire [190:0] _GEN_382; // @[pageswappergcm.scala 880:5:@6082.12]
  wire [2:0] _GEN_383; // @[pageswappergcm.scala 880:5:@6082.12]
  wire [127:0] _GEN_384; // @[pageswappergcm.scala 880:5:@6082.12]
  wire [31:0] _GEN_385; // @[pageswappergcm.scala 880:5:@6082.12]
  wire [190:0] _GEN_386; // @[pageswappergcm.scala 873:5:@6074.10]
  wire [2:0] _GEN_387; // @[pageswappergcm.scala 873:5:@6074.10]
  wire [127:0] _GEN_388; // @[pageswappergcm.scala 873:5:@6074.10]
  wire [31:0] _GEN_389; // @[pageswappergcm.scala 873:5:@6074.10]
  wire [63:0] _GEN_390; // @[pageswappergcm.scala 866:5:@6066.8]
  wire [2:0] _GEN_391; // @[pageswappergcm.scala 866:5:@6066.8]
  wire [190:0] _GEN_392; // @[pageswappergcm.scala 866:5:@6066.8]
  wire [127:0] _GEN_393; // @[pageswappergcm.scala 866:5:@6066.8]
  wire [31:0] _GEN_394; // @[pageswappergcm.scala 866:5:@6066.8]
  wire [2:0] _GEN_395; // @[pageswappergcm.scala 863:5:@6061.6]
  wire [63:0] _GEN_396; // @[pageswappergcm.scala 863:5:@6061.6]
  wire [190:0] _GEN_397; // @[pageswappergcm.scala 863:5:@6061.6]
  wire [127:0] _GEN_398; // @[pageswappergcm.scala 863:5:@6061.6]
  wire [31:0] _GEN_399; // @[pageswappergcm.scala 863:5:@6061.6]
  wire [38:0] _GEN_400; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_401; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [1:0] _GEN_402; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_403; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [1:0] _GEN_404; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_409; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_410; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_411; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_412; // @[pageswappergcm.scala 576:3:@5795.4]
  wire  _GEN_413; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_414; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [2:0] poStateNext; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_416; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_417; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_418; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_419; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [31:0] _GEN_420; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [2:0] _GEN_421; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [63:0] _GEN_422; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [190:0] _GEN_423; // @[pageswappergcm.scala 576:3:@5795.4]
  wire [127:0] _GEN_424; // @[pageswappergcm.scala 576:3:@5795.4]
  randomgen rndgenm ( // @[pageswappergcm.scala 28:23:@5256.4]
    .clock(rndgenm_clock),
    .reset(rndgenm_reset),
    .io_out(rndgenm_io_out),
    .io_en(rndgenm_io_en),
    .io_done(rndgenm_io_done)
  );
  counter cntrm ( // @[pageswappergcm.scala 29:23:@5259.4]
    .clock(cntrm_clock),
    .io_get(cntrm_io_get),
    .io_out(cntrm_io_out),
    .io_reset(cntrm_io_reset),
    .io_init(cntrm_io_init)
  );
  ivFileMac vfm ( // @[pageswappergcm.scala 30:23:@5262.4]
    .clock(vfm_clock),
    .reset(vfm_reset),
    .io_rdata(vfm_io_rdata),
    .io_wdata(vfm_io_wdata),
    .io_addr(vfm_io_addr),
    .io_cmd(vfm_io_cmd)
  );
  aesctr aesm ( // @[pageswappergcm.scala 31:23:@5265.4]
    .clock(aesm_clock),
    .reset(aesm_reset),
    .io_intVect(aesm_io_intVect),
    .io_newR(aesm_io_newR),
    .io_out(aesm_io_out),
    .io_data(aesm_io_data),
    .io_en(aesm_io_en),
    .io_key(aesm_io_key)
  );
  g128Multiplay gmultm ( // @[pageswappergcm.scala 33:22:@5268.4]
    .io_x(gmultm_io_x),
    .io_y(gmultm_io_y),
    .io_out(gmultm_io_out)
  );
  assign start = ConfReg_0[0]; // @[pageswappergcm.scala 125:25:@5337.4]
  assign currOperation = ConfReg_0[3:1]; // @[pageswappergcm.scala 126:33:@5338.4]
  assign aesDone = ConfReg_9[2]; // @[pageswappergcm.scala 128:27:@5339.4]
  assign _T_216 = {ConfReg_1,ConfReg_0}; // @[Cat.scala 30:58:@5340.4]
  assign _T_217 = {ConfReg_3,ConfReg_2}; // @[Cat.scala 30:58:@5341.4]
  assign aesdecInput = {_T_217,_T_216}; // @[Cat.scala 30:58:@5342.4]
  assign _T_219 = currOperation == 3'h1; // @[pageswappergcm.scala 130:37:@5343.4]
  assign _T_221 = currOperation == 3'h3; // @[pageswappergcm.scala 130:63:@5344.4]
  assign _T_222 = _T_219 | _T_221; // @[pageswappergcm.scala 130:46:@5345.4]
  assign _T_223 = {ConfReg_11,ConfReg_10}; // @[Cat.scala 30:58:@5346.4]
  assign _T_224 = {ConfReg_13,ConfReg_12}; // @[Cat.scala 30:58:@5347.4]
  assign _T_225 = {_T_224,_T_223}; // @[Cat.scala 30:58:@5348.4]
  assign aesInOut = _T_222 ? aesdecInput : _T_225; // @[pageswappergcm.scala 130:21:@5349.4]
  assign moduleReady = ConfReg_9[1]; // @[pageswappergcm.scala 134:31:@5350.4]
  assign _T_238 = aesInOut ^ tag; // @[pageswappergcm.scala 145:82:@5358.4]
  assign _T_239 = aesdecInput ^ tag; // @[pageswappergcm.scala 145:102:@5359.4]
  assign _T_240 = _T_222 ? _T_238 : _T_239; // @[pageswappergcm.scala 145:24:@5360.4]
  assign _T_241 = aesDone ? _T_240 : tag; // @[pageswappergcm.scala 144:20:@5361.4]
  assign _GEN_425 = {{7'd0}, ConfReg_2}; // @[pageswappergcm.scala 147:31:@5362.4]
  assign _T_242 = _GEN_425 << 7; // @[pageswappergcm.scala 147:31:@5362.4]
  assign _GEN_426 = {{89'd0}, _T_242}; // @[pageswappergcm.scala 147:37:@5363.4]
  assign _T_243 = _GEN_426 ^ tag; // @[pageswappergcm.scala 147:37:@5363.4]
  assign _T_244 = 2'h3 == tagState; // @[Mux.scala 46:19:@5364.4]
  assign _T_245 = _T_244 ? _T_243 : 128'h0; // @[Mux.scala 46:16:@5365.4]
  assign _T_246 = 2'h2 == tagState; // @[Mux.scala 46:19:@5366.4]
  assign _T_247 = _T_246 ? _T_241 : _T_245; // @[Mux.scala 46:16:@5367.4]
  assign _T_248 = 2'h1 == tagState; // @[Mux.scala 46:19:@5368.4]
  assign _T_249 = _T_248 ? 128'h0 : _T_247; // @[Mux.scala 46:16:@5369.4]
  assign _T_251 = moduleReady == 1'h0; // @[pageswappergcm.scala 151:28:@5371.4]
  assign _T_253 = tagState == 2'h1; // @[pageswappergcm.scala 151:53:@5372.4]
  assign _T_255 = aesDone ? aesInOut : 128'h0; // @[pageswappergcm.scala 151:64:@5373.4]
  assign _T_256 = _T_253 ? _T_255 : IVTag; // @[pageswappergcm.scala 151:43:@5374.4]
  assign _T_257 = _T_251 ? 128'h0 : _T_256; // @[pageswappergcm.scala 151:15:@5375.4]
  assign _T_260 = aesDone & tagUp; // @[pageswappergcm.scala 155:27:@5378.4]
  assign _T_261 = _T_260 ? gmultm_io_out : tag; // @[pageswappergcm.scala 155:18:@5379.4]
  assign _T_263 = cleanupState == 2'h0; // @[pageswappergcm.scala 156:33:@5380.4]
  assign _T_264 = gmultm_io_out ^ IVTag; // @[pageswappergcm.scala 156:71:@5381.4]
  assign _T_265 = _T_263 ? gmultm_io_out : _T_264; // @[pageswappergcm.scala 156:19:@5382.4]
  assign _T_267 = _T_244 ? _T_265 : tag; // @[Mux.scala 46:16:@5384.4]
  assign _T_269 = _T_246 ? _T_261 : _T_267; // @[Mux.scala 46:16:@5386.4]
  assign _T_270 = initState != 3'h6; // @[pageswappergcm.scala 160:31:@5388.4]
  assign _T_274 = initState == 3'h4; // @[pageswappergcm.scala 173:56:@5392.4]
  assign _T_275 = _T_251 & _T_274; // @[pageswappergcm.scala 173:43:@5393.4]
  assign _T_279 = _T_274 & _T_251; // @[pageswappergcm.scala 175:48:@5398.4]
  assign _T_281 = _T_279 ? rndgenm_io_out : 64'h0; // @[pageswappergcm.scala 175:23:@5399.4]
  assign cond1 = poState == 3'h0; // @[pageswappergcm.scala 177:24:@5401.4]
  assign cond2 = blockCounter < ConfReg_2; // @[pageswappergcm.scala 178:28:@5402.4]
  assign _T_283 = poState == 3'h1; // @[pageswappergcm.scala 180:35:@5404.4]
  assign _T_284 = _T_283 & cond2; // @[pageswappergcm.scala 180:48:@5405.4]
  assign _T_285 = cond1 | _T_284; // @[pageswappergcm.scala 180:22:@5406.4]
  assign cond4 = _T_285 & start; // @[pageswappergcm.scala 180:60:@5407.4]
  assign _T_287 = _T_283 & io_memio_ready; // @[pageswappergcm.scala 181:48:@5409.4]
  assign _T_288 = _T_287 & cond2; // @[pageswappergcm.scala 181:66:@5410.4]
  assign _T_289 = cond1 | _T_288; // @[pageswappergcm.scala 181:22:@5411.4]
  assign cond5 = _T_289 & start; // @[pageswappergcm.scala 181:78:@5412.4]
  assign _T_290 = poState == 3'h6; // @[pageswappergcm.scala 183:26:@5413.4]
  assign _T_291 = aesm_io_newR & cond2; // @[pageswappergcm.scala 183:53:@5414.4]
  assign _T_292 = _T_290 | _T_291; // @[pageswappergcm.scala 183:37:@5415.4]
  assign newc24 = _T_292 & start; // @[pageswappergcm.scala 183:64:@5416.4]
  assign _T_298 = 3'h4 == currOperation; // @[Mux.scala 46:19:@5417.4]
  assign _T_299 = _T_298 ? newc24 : 1'h0; // @[Mux.scala 46:16:@5418.4]
  assign _T_300 = 3'h2 == currOperation; // @[Mux.scala 46:19:@5419.4]
  assign _T_301 = _T_300 ? newc24 : _T_299; // @[Mux.scala 46:16:@5420.4]
  assign _T_302 = 3'h3 == currOperation; // @[Mux.scala 46:19:@5421.4]
  assign _T_303 = _T_302 ? cond4 : _T_301; // @[Mux.scala 46:16:@5422.4]
  assign _T_304 = 3'h1 == currOperation; // @[Mux.scala 46:19:@5423.4]
  assign cond = _T_304 ? cond5 : _T_303; // @[Mux.scala 46:16:@5424.4]
  assign newC = _T_251 ? 1'h0 : cond; // @[pageswappergcm.scala 192:14:@5426.4]
  assign _T_311 = cleanupState == 2'h2; // @[pageswappergcm.scala 206:44:@5428.4]
  assign _T_314 = _T_311 ? 2'h2 : 2'h0; // @[pageswappergcm.scala 206:30:@5429.4]
  assign _T_316 = 3'h0 == poState; // @[Mux.scala 46:19:@5430.4]
  assign _T_317 = _T_316 ? 3'h6 : 3'h0; // @[Mux.scala 46:16:@5431.4]
  assign _T_318 = 3'h5 == poState; // @[Mux.scala 46:19:@5432.4]
  assign x1 = _T_318 ? {{1'd0}, _T_314} : _T_317; // @[Mux.scala 46:16:@5433.4]
  assign _T_325 = 2'h2 == cleanupState; // @[Mux.scala 46:19:@5434.4]
  assign _T_326 = _T_325 ? 2'h2 : 2'h0; // @[Mux.scala 46:16:@5435.4]
  assign _T_327 = 2'h0 == cleanupState; // @[Mux.scala 46:19:@5436.4]
  assign _T_328 = _T_327 ? 3'h5 : {{1'd0}, _T_326}; // @[Mux.scala 46:16:@5437.4]
  assign _T_330 = 3'h1 == poState; // @[Mux.scala 46:19:@5438.4]
  assign x3 = _T_318 ? _T_328 : {{2'd0}, _T_330}; // @[Mux.scala 46:16:@5441.4]
  assign _T_341 = _T_318 ? 2'h3 : 2'h0; // @[Mux.scala 46:16:@5445.4]
  assign _T_342 = 3'h6 == poState; // @[Mux.scala 46:19:@5446.4]
  assign x2 = _T_342 ? {{1'd0}, start} : _T_341; // @[Mux.scala 46:16:@5447.4]
  assign _T_350 = blockCounter > 32'h1; // @[pageswappergcm.scala 231:47:@5450.4]
  assign _T_353 = _T_350 ? 2'h2 : 2'h0; // @[pageswappergcm.scala 231:32:@5451.4]
  assign _T_355 = blockCounter == 32'h0; // @[pageswappergcm.scala 232:43:@5452.4]
  assign _T_358 = _T_355 ? 2'h3 : 2'h0; // @[pageswappergcm.scala 232:29:@5453.4]
  assign _T_359 = 3'h2 == poState; // @[Mux.scala 46:19:@5454.4]
  assign _T_360 = _T_359 ? _T_358 : 2'h0; // @[Mux.scala 46:16:@5455.4]
  assign _T_361 = 3'h3 == poState; // @[Mux.scala 46:19:@5456.4]
  assign _T_362 = _T_361 ? _T_353 : _T_360; // @[Mux.scala 46:16:@5457.4]
  assign x4 = _T_342 ? {{1'd0}, start} : _T_362; // @[Mux.scala 46:16:@5459.4]
  assign _T_370 = _T_298 ? x4 : 2'h0; // @[Mux.scala 46:16:@5461.4]
  assign _T_372 = _T_302 ? x3 : {{1'd0}, _T_370}; // @[Mux.scala 46:16:@5463.4]
  assign _T_374 = _T_300 ? {{1'd0}, x2} : _T_372; // @[Mux.scala 46:16:@5465.4]
  assign _T_376 = _T_304 ? x1 : _T_374; // @[Mux.scala 46:16:@5467.4]
  assign _T_378 = poState == 3'h5; // @[pageswappergcm.scala 250:27:@5469.4]
  assign _T_380 = _T_378 ? 32'h0 : ConfReg_3; // @[pageswappergcm.scala 250:18:@5470.4]
  assign _T_386 = blockCounter - 32'h2; // @[pageswappergcm.scala 254:70:@5472.4]
  assign _T_387 = $unsigned(_T_386); // @[pageswappergcm.scala 254:70:@5473.4]
  assign _T_388 = _T_387[31:0]; // @[pageswappergcm.scala 254:70:@5474.4]
  assign _T_389 = _T_350 ? _T_388 : blockCounter; // @[pageswappergcm.scala 254:35:@5475.4]
  assign _T_391 = _T_361 ? _T_389 : 32'h0; // @[Mux.scala 46:16:@5477.4]
  assign _T_393 = _T_298 ? _T_391 : ConfReg_3; // @[Mux.scala 46:16:@5479.4]
  assign _T_395 = _T_302 ? _T_380 : _T_393; // @[Mux.scala 46:16:@5481.4]
  assign _GEN_427 = {{255'd0}, sessionIv}; // @[pageswappergcm.scala 264:40:@5483.4]
  assign _T_400 = _GEN_427 << 8'h80; // @[pageswappergcm.scala 264:40:@5483.4]
  assign _GEN_428 = {{255'd0}, tag}; // @[pageswappergcm.scala 264:49:@5484.4]
  assign _T_401 = _T_400 | _GEN_428; // @[pageswappergcm.scala 264:49:@5484.4]
  assign _T_402 = {1'h1,_T_401}; // @[Cat.scala 30:58:@5485.4]
  assign _T_408 = {1'h0,_T_401}; // @[Cat.scala 30:58:@5488.4]
  assign _GEN_433 = {{255'd0}, aesInOut}; // @[pageswappergcm.scala 267:39:@5492.4]
  assign _T_418 = _GEN_433 << 8'h80; // @[pageswappergcm.scala 267:39:@5492.4]
  assign _T_419 = _T_418 | _GEN_433; // @[pageswappergcm.scala 267:48:@5493.4]
  assign _T_420 = {1'h1,_T_419}; // @[Cat.scala 30:58:@5494.4]
  assign _T_422 = _T_298 ? _T_420 : 384'h0; // @[Mux.scala 46:16:@5496.4]
  assign _T_424 = _T_302 ? _T_402 : _T_422; // @[Mux.scala 46:16:@5498.4]
  assign _T_426 = _T_300 ? _T_408 : _T_424; // @[Mux.scala 46:16:@5500.4]
  assign _T_428 = _T_304 ? _T_402 : _T_426; // @[Mux.scala 46:16:@5502.4]
  assign _GEN_435 = {{127'd0}, nonce}; // @[pageswappergcm.scala 277:30:@5504.4]
  assign _T_430 = _GEN_435 << 7'h40; // @[pageswappergcm.scala 277:30:@5504.4]
  assign _GEN_436 = {{127'd0}, cntrm_io_out}; // @[pageswappergcm.scala 277:38:@5505.4]
  assign _T_431 = _T_430 | _GEN_436; // @[pageswappergcm.scala 277:38:@5505.4]
  assign cv13 = newC ? _T_431 : {{63'd0}, curriv}; // @[pageswappergcm.scala 277:17:@5506.4]
  assign _T_435 = cond1 & _T_355; // @[pageswappergcm.scala 278:37:@5509.4]
  assign _T_436 = poState == 3'h3; // @[pageswappergcm.scala 279:18:@5510.4]
  assign _T_438 = curriv + 128'h1; // @[pageswappergcm.scala 279:40:@5511.4]
  assign _T_439 = _T_438[127:0]; // @[pageswappergcm.scala 279:40:@5512.4]
  assign _T_440 = _T_436 ? _T_439 : curriv; // @[pageswappergcm.scala 279:8:@5513.4]
  assign cv2 = _T_435 ? vfm_io_rdata : _T_440; // @[pageswappergcm.scala 278:17:@5514.4]
  assign _T_446 = _T_298 ? cv2 : curriv; // @[Mux.scala 46:16:@5516.4]
  assign _T_448 = _T_300 ? cv2 : _T_446; // @[Mux.scala 46:16:@5518.4]
  assign _T_450 = _T_302 ? cv13 : {{63'd0}, _T_448}; // @[Mux.scala 46:16:@5520.4]
  assign xcv = _T_304 ? cv13 : _T_450; // @[Mux.scala 46:16:@5522.4]
  assign _T_454 = cond1 ? xcv : {{63'd0}, sessionIv}; // @[pageswappergcm.scala 298:20:@5525.4]
  assign _T_460 = _T_378 ? vfm_io_rdata : sessionIv; // @[pageswappergcm.scala 300:20:@5529.4]
  assign _T_462 = poState == 3'h2; // @[pageswappergcm.scala 301:30:@5530.4]
  assign _T_465 = _T_462 & _T_355; // @[pageswappergcm.scala 301:41:@5532.4]
  assign _T_466 = _T_465 ? vfm_io_rdata : sessionIv; // @[pageswappergcm.scala 301:20:@5533.4]
  assign _T_468 = _T_298 ? _T_466 : sessionIv; // @[Mux.scala 46:16:@5535.4]
  assign _T_470 = _T_300 ? _T_460 : _T_468; // @[Mux.scala 46:16:@5537.4]
  assign _T_472 = _T_302 ? _T_454 : {{63'd0}, _T_470}; // @[Mux.scala 46:16:@5539.4]
  assign _T_474 = _T_304 ? _T_454 : _T_472; // @[Mux.scala 46:16:@5541.4]
  assign _T_476 = blockCounter < 32'h1; // @[pageswappergcm.scala 313:31:@5543.4]
  assign bcg1 = _T_476 ? 1'h0 : aesDone; // @[pageswappergcm.scala 313:17:@5545.4]
  assign _T_480 = blockCounter <= 32'h1; // @[pageswappergcm.scala 314:31:@5546.4]
  assign bcg2 = _T_480 ? 1'h0 : aesDone; // @[pageswappergcm.scala 314:17:@5548.4]
  assign _T_489 = _T_298 ? bcg2 : 1'h0; // @[Mux.scala 46:16:@5550.4]
  assign _T_491 = _T_302 ? bcg1 : _T_489; // @[Mux.scala 46:16:@5552.4]
  assign _T_493 = _T_300 ? bcg2 : _T_491; // @[Mux.scala 46:16:@5554.4]
  assign _T_495 = _T_304 ? bcg1 : _T_493; // @[Mux.scala 46:16:@5556.4]
  assign _T_497 = ConfReg_4 != 32'h0; // @[pageswappergcm.scala 340:24:@5558.4]
  assign _T_498 = ConfReg_9[4]; // @[pageswappergcm.scala 341:28:@5560.4]
  assign _T_503 = _T_283 ? io_memio_rdata : currBlockBuff; // @[pageswappergcm.scala 346:43:@5564.4]
  assign _T_504 = _T_253 ? 128'h0 : _T_503; // @[pageswappergcm.scala 346:18:@5565.4]
  assign _T_508 = _T_253 ? 128'h0 : vfm_io_rdata; // @[pageswappergcm.scala 347:18:@5567.4]
  assign _T_512 = _T_298 ? aesdecInput : currBlockBuff; // @[Mux.scala 46:16:@5569.4]
  assign _T_514 = _T_300 ? aesdecInput : _T_512; // @[Mux.scala 46:16:@5571.4]
  assign _T_516 = _T_302 ? _T_508 : _T_514; // @[Mux.scala 46:16:@5573.4]
  assign cb = _T_304 ? _T_504 : _T_516; // @[Mux.scala 46:16:@5575.4]
  assign _T_522 = initState == 3'h5; // @[pageswappergcm.scala 357:46:@5580.4]
  assign _T_524 = _T_251 ? _T_522 : _T_462; // @[pageswappergcm.scala 357:14:@5582.4]
  assign _T_528 = _T_251 ? 128'h0 : curriv; // @[pageswappergcm.scala 359:25:@5586.4]
  assign _T_533 = _T_251 ? 128'h0 : cb; // @[pageswappergcm.scala 363:29:@5589.4]
  assign _T_543 = _T_355 ? 128'h0 : cb; // @[pageswappergcm.scala 365:29:@5593.4]
  assign _T_550 = _T_298 ? _T_543 : cb; // @[Mux.scala 46:16:@5597.4]
  assign _T_552 = _T_300 ? _T_543 : _T_550; // @[Mux.scala 46:16:@5599.4]
  assign _T_554 = _T_302 ? _T_533 : _T_552; // @[Mux.scala 46:16:@5601.4]
  assign _T_556 = _T_304 ? _T_533 : _T_554; // @[Mux.scala 46:16:@5603.4]
  assign socmselect = io_mainMemio_addr < 14'h2000; // @[pageswappergcm.scala 387:38:@5622.4]
  assign _T_583 = io_mainMemio_addr >= 14'h2000; // @[pageswappergcm.scala 388:44:@5623.4]
  assign _T_586 = 14'h2000 + 14'h9; // @[pageswappergcm.scala 388:123:@5624.4]
  assign _T_587 = _T_586[13:0]; // @[pageswappergcm.scala 388:123:@5625.4]
  assign _T_588 = io_mainMemio_addr <= _T_587; // @[pageswappergcm.scala 388:94:@5626.4]
  assign validConfAddress = _T_583 & _T_588; // @[pageswappergcm.scala 388:73:@5627.4]
  assign _T_590 = currOperation == 3'h5; // @[pageswappergcm.scala 393:45:@5630.4]
  assign _T_591 = _T_590 & socmselect; // @[pageswappergcm.scala 393:54:@5631.4]
  assign _T_598 = _T_591 ? io_mainMemio_we : 1'h0; // @[pageswappergcm.scala 394:29:@5636.4]
  assign _T_603 = _T_591 ? io_mainMemio_en : 1'h0; // @[pageswappergcm.scala 395:29:@5640.4]
  assign confaddr = io_mainMemio_addr[3:0]; // @[pageswappergcm.scala 398:35:@5642.4]
  assign _T_811 = aesm_io_out[63:32]; // @[pageswappergcm.scala 635:42:@5848.20]
  assign _GEN_121 = aesm_io_newR ? _T_811 : ConfReg_1; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_158 = _T_462 ? _GEN_121 : ConfReg_1; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_175 = _T_283 ? ConfReg_1 : _GEN_158; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_191 = cond1 ? ConfReg_1 : _GEN_175; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_206 = _T_290 ? ConfReg_1 : _GEN_191; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_330 = _T_222 ? _GEN_206 : ConfReg_1; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_351 = start ? _GEN_330 : ConfReg_1; // @[pageswappergcm.scala 580:5:@5797.6]
  assign ConfRegWire_1 = moduleReady ? _GEN_351 : ConfReg_1; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _T_810 = aesm_io_out[31:0]; // @[pageswappergcm.scala 634:42:@5846.20]
  assign _GEN_120 = aesm_io_newR ? _T_810 : ConfReg_0; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_157 = _T_462 ? _GEN_120 : ConfReg_0; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_174 = _T_283 ? ConfReg_0 : _GEN_157; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_190 = cond1 ? ConfReg_0 : _GEN_174; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_205 = _T_290 ? ConfReg_0 : _GEN_190; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_329 = _T_222 ? _GEN_205 : ConfReg_0; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_350 = start ? _GEN_329 : ConfReg_0; // @[pageswappergcm.scala 580:5:@5797.6]
  assign ConfRegWire_0 = moduleReady ? _GEN_350 : ConfReg_0; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_4 = 4'h1 == confaddr ? ConfRegWire_1 : ConfRegWire_0; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _T_812 = aesm_io_out[95:64]; // @[pageswappergcm.scala 636:42:@5850.20]
  assign _GEN_122 = aesm_io_newR ? _T_812 : ConfReg_2; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_159 = _T_462 ? _GEN_122 : ConfReg_2; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_176 = _T_283 ? ConfReg_2 : _GEN_159; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_192 = cond1 ? ConfReg_2 : _GEN_176; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_207 = _T_290 ? ConfReg_2 : _GEN_192; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_331 = _T_222 ? _GEN_207 : ConfReg_2; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_352 = start ? _GEN_331 : ConfReg_2; // @[pageswappergcm.scala 580:5:@5797.6]
  assign ConfRegWire_2 = moduleReady ? _GEN_352 : ConfReg_2; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_5 = 4'h2 == confaddr ? ConfRegWire_2 : _GEN_4; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _T_813 = aesm_io_out[127:96]; // @[pageswappergcm.scala 637:42:@5852.20]
  assign _GEN_123 = aesm_io_newR ? _T_813 : ConfReg_3; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_160 = _T_462 ? _GEN_123 : ConfReg_3; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_177 = _T_283 ? ConfReg_3 : _GEN_160; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_193 = cond1 ? ConfReg_3 : _GEN_177; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_208 = _T_290 ? ConfReg_3 : _GEN_193; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_332 = _T_222 ? _GEN_208 : ConfReg_3; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_353 = start ? _GEN_332 : ConfReg_3; // @[pageswappergcm.scala 580:5:@5797.6]
  assign ConfRegWire_3 = moduleReady ? _GEN_353 : ConfReg_3; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_6 = 4'h3 == confaddr ? ConfRegWire_3 : _GEN_5; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_7 = 4'h4 == confaddr ? ConfReg_4 : _GEN_6; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_8 = 4'h5 == confaddr ? ConfReg_5 : _GEN_7; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_9 = 4'h6 == confaddr ? ConfReg_6 : _GEN_8; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_10 = 4'h7 == confaddr ? ConfReg_7 : _GEN_9; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_11 = 4'h8 == confaddr ? ConfReg_8 : _GEN_10; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_12 = 4'h9 == confaddr ? ConfReg_9 : _GEN_11; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_13 = 4'ha == confaddr ? ConfReg_10 : _GEN_12; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_14 = 4'hb == confaddr ? ConfReg_11 : _GEN_13; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_15 = 4'hc == confaddr ? ConfReg_12 : _GEN_14; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _GEN_16 = 4'hd == confaddr ? ConfReg_13 : _GEN_15; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _T_608 = _T_591 ? io_socMemio_rdata : _GEN_16; // @[pageswappergcm.scala 412:29:@5645.4]
  assign _T_611 = io_mainMemio_en & io_mainMemio_valid; // @[pageswappergcm.scala 416:55:@5647.4]
  assign _T_616 = _T_590 ? io_socMemio_ready : 1'h0; // @[pageswappergcm.scala 417:41:@5649.4]
  assign _T_618 = socmselect ? _T_616 : 1'h0; // @[Mux.scala 46:16:@5651.4]
  assign _T_619 = 1'h0 == socmselect; // @[Mux.scala 46:19:@5652.4]
  assign _T_620 = _T_619 ? _T_611 : _T_618; // @[Mux.scala 46:16:@5653.4]
  assign _T_625 = 4'h9 == confaddr; // @[Mux.scala 46:19:@5656.4]
  assign confMask = _T_625 ? 32'h1f : 32'h0; // @[Mux.scala 46:16:@5657.4]
  assign _T_627 = currOperation == 3'h2; // @[pageswappergcm.scala 437:42:@5658.4]
  assign _T_629 = currOperation == 3'h4; // @[pageswappergcm.scala 437:69:@5659.4]
  assign _T_630 = _T_627 | _T_629; // @[pageswappergcm.scala 437:51:@5660.4]
  assign _T_631 = ConfReg_9[5]; // @[pageswappergcm.scala 437:90:@5661.4]
  assign pindataReady = _T_630 ? _T_631 : 1'h0; // @[pageswappergcm.scala 437:25:@5662.4]
  assign _T_638 = ConfReg_9[6]; // @[pageswappergcm.scala 438:91:@5666.4]
  assign poutdataReady = _T_222 ? _T_638 : 1'h0; // @[pageswappergcm.scala 438:26:@5667.4]
  assign _T_641 = ~ socmselect; // @[pageswappergcm.scala 447:14:@5671.6]
  assign _T_642 = _T_641 & validConfAddress; // @[pageswappergcm.scala 447:26:@5672.6]
  assign _T_643 = ~ confMask; // @[pageswappergcm.scala 451:48:@5675.10]
  assign _T_644 = io_mainMemio_wdata & _T_643; // @[pageswappergcm.scala 451:45:@5676.10]
  assign _T_646 = confMask == 32'h0; // @[pageswappergcm.scala 455:35:@5677.10]
  assign _T_647 = ~ _T_646; // @[pageswappergcm.scala 456:19:@5678.10]
  assign _GEN_17 = 4'h1 == confaddr ? ConfReg_1 : ConfReg_0; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_18 = 4'h2 == confaddr ? ConfReg_2 : _GEN_17; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_19 = 4'h3 == confaddr ? ConfReg_3 : _GEN_18; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_20 = 4'h4 == confaddr ? ConfReg_4 : _GEN_19; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_21 = 4'h5 == confaddr ? ConfReg_5 : _GEN_20; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_22 = 4'h6 == confaddr ? ConfReg_6 : _GEN_21; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_23 = 4'h7 == confaddr ? ConfReg_7 : _GEN_22; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_24 = 4'h8 == confaddr ? ConfReg_8 : _GEN_23; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_25 = 4'h9 == confaddr ? ConfReg_9 : _GEN_24; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_26 = 4'ha == confaddr ? ConfReg_10 : _GEN_25; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_27 = 4'hb == confaddr ? ConfReg_11 : _GEN_26; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_28 = 4'hc == confaddr ? ConfReg_12 : _GEN_27; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_29 = 4'hd == confaddr ? ConfReg_13 : _GEN_28; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _T_656 = _GEN_29 | _T_644; // @[pageswappergcm.scala 463:85:@5682.12]
  assign _GEN_30 = 4'h0 == confaddr ? _T_656 : ConfReg_0; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_31 = 4'h1 == confaddr ? _T_656 : ConfReg_1; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_32 = 4'h2 == confaddr ? _T_656 : ConfReg_2; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_35 = 4'h5 == confaddr ? _T_656 : ConfReg_5; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_36 = 4'h6 == confaddr ? _T_656 : ConfReg_6; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_37 = 4'h7 == confaddr ? _T_656 : ConfReg_7; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_38 = 4'h8 == confaddr ? _T_656 : ConfReg_8; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_39 = 4'h9 == confaddr ? _T_656 : ConfReg_9; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_40 = 4'ha == confaddr ? _T_656 : ConfReg_10; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_41 = 4'hb == confaddr ? _T_656 : ConfReg_11; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_42 = 4'hc == confaddr ? _T_656 : ConfReg_12; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_43 = 4'hd == confaddr ? _T_656 : ConfReg_13; // @[pageswappergcm.scala 463:50:@5683.12]
  assign _GEN_44 = 4'h0 == confaddr ? _T_644 : ConfReg_0; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_45 = 4'h1 == confaddr ? _T_644 : ConfReg_1; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_46 = 4'h2 == confaddr ? _T_644 : ConfReg_2; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_49 = 4'h5 == confaddr ? _T_644 : ConfReg_5; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_50 = 4'h6 == confaddr ? _T_644 : ConfReg_6; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_51 = 4'h7 == confaddr ? _T_644 : ConfReg_7; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_52 = 4'h8 == confaddr ? _T_644 : ConfReg_8; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_53 = 4'h9 == confaddr ? _T_644 : ConfReg_9; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_54 = 4'ha == confaddr ? _T_644 : ConfReg_10; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_55 = 4'hb == confaddr ? _T_644 : ConfReg_11; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_56 = 4'hc == confaddr ? _T_644 : ConfReg_12; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_57 = 4'hd == confaddr ? _T_644 : ConfReg_13; // @[pageswappergcm.scala 472:50:@5687.12]
  assign _GEN_58 = _T_647 ? _GEN_30 : _GEN_44; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_59 = _T_647 ? _GEN_31 : _GEN_45; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_60 = _T_647 ? _GEN_32 : _GEN_46; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_63 = _T_647 ? _GEN_35 : _GEN_49; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_64 = _T_647 ? _GEN_36 : _GEN_50; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_65 = _T_647 ? _GEN_37 : _GEN_51; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_66 = _T_647 ? _GEN_38 : _GEN_52; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_67 = _T_647 ? _GEN_39 : _GEN_53; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_68 = _T_647 ? _GEN_40 : _GEN_54; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_69 = _T_647 ? _GEN_41 : _GEN_55; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_70 = _T_647 ? _GEN_42 : _GEN_56; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _GEN_71 = _T_647 ? _GEN_43 : _GEN_57; // @[pageswappergcm.scala 457:14:@5679.10]
  assign _T_667 = currOperation == 3'h0; // @[pageswappergcm.scala 476:95:@5692.10]
  assign _T_668 = _T_630 | _T_667; // @[pageswappergcm.scala 476:77:@5693.10]
  assign _T_671 = confaddr == 4'h8; // @[pageswappergcm.scala 476:132:@5695.10]
  assign _T_672 = _T_668 & _T_671; // @[pageswappergcm.scala 476:105:@5696.10]
  assign _T_675 = 8'h1 << 3'h5; // @[pageswappergcm.scala 479:47:@5698.12]
  assign _GEN_437 = {{24'd0}, _T_675}; // @[pageswappergcm.scala 479:41:@5699.12]
  assign _T_676 = ConfReg_9 | _GEN_437; // @[pageswappergcm.scala 479:41:@5699.12]
  assign _GEN_72 = _T_672 ? _T_676 : _GEN_67; // @[pageswappergcm.scala 478:14:@5697.10]
  assign _GEN_73 = io_mainMemio_we ? _GEN_58 : ConfReg_0; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_74 = io_mainMemio_we ? _GEN_59 : ConfReg_1; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_75 = io_mainMemio_we ? _GEN_60 : ConfReg_2; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_78 = io_mainMemio_we ? _GEN_63 : ConfReg_5; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_79 = io_mainMemio_we ? _GEN_64 : ConfReg_6; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_80 = io_mainMemio_we ? _GEN_65 : ConfReg_7; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_81 = io_mainMemio_we ? _GEN_66 : ConfReg_8; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_82 = io_mainMemio_we ? _GEN_72 : ConfReg_9; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_83 = io_mainMemio_we ? _GEN_68 : ConfReg_10; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_84 = io_mainMemio_we ? _GEN_69 : ConfReg_11; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_85 = io_mainMemio_we ? _GEN_70 : ConfReg_12; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_86 = io_mainMemio_we ? _GEN_71 : ConfReg_13; // @[pageswappergcm.scala 450:12:@5674.8]
  assign _GEN_87 = _T_642 ? _GEN_73 : ConfReg_0; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_88 = _T_642 ? _GEN_74 : ConfReg_1; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_89 = _T_642 ? _GEN_75 : ConfReg_2; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_92 = _T_642 ? _GEN_78 : ConfReg_5; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_93 = _T_642 ? _GEN_79 : ConfReg_6; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_94 = _T_642 ? _GEN_80 : ConfReg_7; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_95 = _T_642 ? _GEN_81 : ConfReg_8; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_96 = _T_642 ? _GEN_82 : ConfReg_9; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_97 = _T_642 ? _GEN_83 : ConfReg_10; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_98 = _T_642 ? _GEN_84 : ConfReg_11; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_99 = _T_642 ? _GEN_85 : ConfReg_12; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_100 = _T_642 ? _GEN_86 : ConfReg_13; // @[pageswappergcm.scala 448:9:@5673.6]
  assign _GEN_101 = _T_611 ? _GEN_87 : ConfReg_0; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_102 = _T_611 ? _GEN_88 : ConfReg_1; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_103 = _T_611 ? _GEN_89 : ConfReg_2; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_106 = _T_611 ? _GEN_92 : ConfReg_5; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_107 = _T_611 ? _GEN_93 : ConfReg_6; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_108 = _T_611 ? _GEN_94 : ConfReg_7; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_109 = _T_611 ? _GEN_95 : ConfReg_8; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_110 = _T_611 ? _GEN_96 : ConfReg_9; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_111 = _T_611 ? _GEN_97 : ConfReg_10; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_112 = _T_611 ? _GEN_98 : ConfReg_11; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_113 = _T_611 ? _GEN_99 : ConfReg_12; // @[pageswappergcm.scala 445:3:@5670.4]
  assign _GEN_114 = _T_611 ? _GEN_100 : ConfReg_13; // @[pageswappergcm.scala 445:3:@5670.4]
  assign vfNotFull = vfm_io_rdata <= 128'hf; // @[pageswappergcm.scala 498:34:@5707.4]
  assign _T_681 = cond1 & vfNotFull; // @[pageswappergcm.scala 502:42:@5709.4]
  assign _T_683 = _T_681 ? vfm_io_rdata : 128'h0; // @[pageswappergcm.scala 502:22:@5710.4]
  assign _T_686 = _T_302 ? blockCounter : 32'h0; // @[Mux.scala 46:16:@5712.4]
  assign conf3 = _T_304 ? _T_683 : {{96'd0}, _T_686}; // @[Mux.scala 46:16:@5714.4]
  assign _T_689 = start ? conf3 : {{96'd0}, ConfReg_3}; // @[pageswappergcm.scala 505:22:@5716.4]
  assign _T_693 = ~ vfNotFull; // @[pageswappergcm.scala 511:44:@5719.4]
  assign _T_694 = cond1 & _T_693; // @[pageswappergcm.scala 511:41:@5720.4]
  assign _T_696 = ConfReg_4 | 32'h1; // @[pageswappergcm.scala 511:68:@5721.4]
  assign _T_697 = _T_694 ? _T_696 : ConfReg_4; // @[pageswappergcm.scala 511:20:@5722.4]
  assign conf4 = _T_304 ? _T_697 : 32'h0; // @[Mux.scala 46:16:@5724.4]
  assign _T_700 = start ? conf4 : ConfReg_4; // @[pageswappergcm.scala 513:22:@5726.4]
  assign _T_713 = _T_300 ? _T_436 : 1'h0; // @[Mux.scala 46:16:@5733.4]
  assign mmenvalid = _T_304 ? _T_283 : _T_713; // @[Mux.scala 46:16:@5735.4]
  assign _T_720 = ConfReg_1[10:0]; // @[pageswappergcm.scala 533:27:@5741.4]
  assign _GEN_438 = {{21'd0}, _T_720}; // @[pageswappergcm.scala 533:63:@5745.4]
  assign _T_725 = _GEN_438 + _T_388; // @[pageswappergcm.scala 533:63:@5745.4]
  assign addr2 = _T_725[31:0]; // @[pageswappergcm.scala 533:63:@5746.4]
  assign _T_727 = _GEN_438 + blockCounter; // @[pageswappergcm.scala 536:63:@5748.4]
  assign addr1 = _T_727[31:0]; // @[pageswappergcm.scala 536:63:@5749.4]
  assign _T_732 = _T_283 ? addr1 : 32'h0; // @[pageswappergcm.scala 541:19:@5751.4]
  assign _T_736 = _T_436 ? addr2 : 32'h0; // @[pageswappergcm.scala 542:19:@5753.4]
  assign _T_738 = _T_300 ? _T_736 : 32'h0; // @[Mux.scala 46:16:@5755.4]
  assign addr = _T_304 ? _T_732 : _T_738; // @[Mux.scala 46:16:@5757.4]
  assign _T_743 = _T_436 & _T_627; // @[pageswappergcm.scala 546:48:@5761.4]
  assign _T_748 = _T_743 ? _T_225 : 128'h0; // @[pageswappergcm.scala 546:25:@5765.4]
  assign nPoState = _T_253 ? 3'h1 : 3'h4; // @[pageswappergcm.scala 552:21:@5769.4]
  assign _T_751 = cond2 ? nPoState : 3'h4; // @[pageswappergcm.scala 559:40:@5770.4]
  assign _T_752 = aesm_io_newR ? _T_751 : 3'h2; // @[pageswappergcm.scala 559:23:@5771.4]
  assign _T_753 = cond2 ? 3'h1 : 3'h5; // @[pageswappergcm.scala 560:47:@5772.4]
  assign _T_754 = poutdataReady ? _T_753 : 3'h4; // @[pageswappergcm.scala 560:29:@5773.4]
  assign _T_757 = io_memio_ready ? 3'h2 : 3'h1; // @[pageswappergcm.scala 561:50:@5775.4]
  assign _T_758 = _T_219 ? _T_757 : 3'h2; // @[pageswappergcm.scala 561:24:@5776.4]
  assign _T_761 = _T_311 ? 3'h6 : 3'h5; // @[pageswappergcm.scala 562:24:@5778.4]
  assign _T_763 = _T_318 ? _T_761 : 3'h6; // @[Mux.scala 46:16:@5780.4]
  assign _T_765 = _T_330 ? _T_758 : _T_763; // @[Mux.scala 46:16:@5782.4]
  assign _T_766 = 3'h4 == poState; // @[Mux.scala 46:19:@5783.4]
  assign _T_767 = _T_766 ? _T_754 : _T_765; // @[Mux.scala 46:16:@5784.4]
  assign _T_769 = _T_359 ? _T_752 : _T_767; // @[Mux.scala 46:16:@5786.4]
  assign _T_771 = _T_316 ? 3'h2 : _T_769; // @[Mux.scala 46:16:@5788.4]
  assign pos13 = _T_342 ? 3'h0 : _T_771; // @[Mux.scala 46:16:@5790.4]
  assign _T_773 = start & moduleReady; // @[pageswappergcm.scala 566:28:@5791.4]
  assign _T_774 = _T_773 ? pos13 : 3'h6; // @[pageswappergcm.scala 566:21:@5792.4]
  assign _T_785 = 35'h1 << 2'h2; // @[pageswappergcm.scala 588:49:@5804.12]
  assign _T_786 = ~ _T_785; // @[pageswappergcm.scala 588:38:@5805.12]
  assign _GEN_440 = {{3'd0}, ConfReg_9}; // @[pageswappergcm.scala 588:36:@5806.12]
  assign _T_787 = _GEN_440 & _T_786; // @[pageswappergcm.scala 588:36:@5806.12]
  assign _GEN_115 = _T_221 ? 32'h20 : _GEN_103; // @[pageswappergcm.scala 595:13:@5813.14]
  assign _GEN_116 = _T_221 ? 2'h0 : cleanupStateNext; // @[pageswappergcm.scala 595:13:@5813.14]
  assign _T_796 = 4'h1 << 2'h2; // @[pageswappergcm.scala 604:46:@5821.16]
  assign _T_797 = ~ _T_796; // @[pageswappergcm.scala 604:41:@5822.16]
  assign _GEN_441 = {{28'd0}, _T_797}; // @[pageswappergcm.scala 604:38:@5823.16]
  assign _T_798 = ConfReg_9 & _GEN_441; // @[pageswappergcm.scala 604:38:@5823.16]
  assign _T_802 = blockCounter + 32'h1; // @[pageswappergcm.scala 616:46:@5828.20]
  assign _T_803 = _T_802[31:0]; // @[pageswappergcm.scala 616:46:@5829.20]
  assign _GEN_117 = io_memio_ready ? _T_803 : blockCounter; // @[pageswappergcm.scala 614:15:@5827.18]
  assign _GEN_118 = _T_221 ? _T_803 : blockCounter; // @[pageswappergcm.scala 621:13:@5835.18]
  assign _GEN_119 = _T_219 ? _GEN_117 : _GEN_118; // @[pageswappergcm.scala 606:13:@5826.16]
  assign _GEN_442 = {{28'd0}, _T_796}; // @[pageswappergcm.scala 655:38:@5864.20]
  assign _T_822 = ConfReg_9 | _GEN_442; // @[pageswappergcm.scala 655:38:@5864.20]
  assign _GEN_124 = aesm_io_newR ? _T_810 : _GEN_106; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_125 = aesm_io_newR ? _T_811 : _GEN_107; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_126 = aesm_io_newR ? _T_812 : _GEN_108; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_127 = aesm_io_newR ? _T_813 : _GEN_109; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_128 = aesm_io_newR ? 1'h1 : tagUp; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _GEN_129 = aesm_io_newR ? _T_822 : _GEN_110; // @[pageswappergcm.scala 632:11:@5845.18]
  assign _T_823 = poState == 3'h4; // @[pageswappergcm.scala 683:28:@5869.18]
  assign _T_827 = 39'h1 << 3'h6; // @[pageswappergcm.scala 691:55:@5873.22]
  assign _T_828 = ~ _T_827; // @[pageswappergcm.scala 691:44:@5874.22]
  assign _GEN_443 = {{7'd0}, ConfReg_9}; // @[pageswappergcm.scala 691:42:@5875.22]
  assign _T_829 = _GEN_443 & _T_828; // @[pageswappergcm.scala 691:42:@5875.22]
  assign _GEN_130 = poutdataReady ? _T_829 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 689:15:@5872.20]
  assign _T_835 = cleanupState == 2'h1; // @[pageswappergcm.scala 708:37:@5888.24]
  assign _T_840 = ConfReg_0 & 32'hfffffffe; // @[pageswappergcm.scala 715:41:@5896.28]
  assign _T_843 = 39'h1 << 3'h4; // @[pageswappergcm.scala 716:53:@5898.28]
  assign _T_844 = _GEN_443 | _T_843; // @[pageswappergcm.scala 716:41:@5899.28]
  assign _GEN_131 = _T_311 ? _T_840 : _GEN_101; // @[pageswappergcm.scala 713:12:@5895.26]
  assign _GEN_132 = _T_311 ? _T_844 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 713:12:@5895.26]
  assign _GEN_133 = _T_311 ? 2'h1 : 2'h3; // @[pageswappergcm.scala 713:12:@5895.26]
  assign _GEN_134 = _T_311 ? 32'h0 : blockCounter; // @[pageswappergcm.scala 713:12:@5895.26]
  assign _GEN_135 = _T_311 ? 2'h0 : cleanupStateNext; // @[pageswappergcm.scala 713:12:@5895.26]
  assign _GEN_136 = _T_835 ? 2'h2 : _GEN_135; // @[pageswappergcm.scala 709:12:@5889.24]
  assign _GEN_137 = _T_835 ? 2'h1 : _GEN_133; // @[pageswappergcm.scala 709:12:@5889.24]
  assign _GEN_138 = _T_835 ? _GEN_101 : _GEN_131; // @[pageswappergcm.scala 709:12:@5889.24]
  assign _GEN_139 = _T_835 ? {{7'd0}, _GEN_110} : _GEN_132; // @[pageswappergcm.scala 709:12:@5889.24]
  assign _GEN_140 = _T_835 ? blockCounter : _GEN_134; // @[pageswappergcm.scala 709:12:@5889.24]
  assign _GEN_141 = _T_263 ? 2'h1 : _GEN_136; // @[pageswappergcm.scala 704:12:@5884.22]
  assign _GEN_142 = _T_263 ? 2'h3 : _GEN_137; // @[pageswappergcm.scala 704:12:@5884.22]
  assign _GEN_143 = _T_263 ? _GEN_101 : _GEN_138; // @[pageswappergcm.scala 704:12:@5884.22]
  assign _GEN_144 = _T_263 ? {{7'd0}, _GEN_110} : _GEN_139; // @[pageswappergcm.scala 704:12:@5884.22]
  assign _GEN_145 = _T_263 ? blockCounter : _GEN_140; // @[pageswappergcm.scala 704:12:@5884.22]
  assign _GEN_146 = _T_378 ? _GEN_142 : tagState; // @[pageswappergcm.scala 697:9:@5881.20]
  assign _GEN_147 = _T_378 ? _GEN_141 : cleanupStateNext; // @[pageswappergcm.scala 697:9:@5881.20]
  assign _GEN_148 = _T_378 ? _GEN_143 : _GEN_101; // @[pageswappergcm.scala 697:9:@5881.20]
  assign _GEN_149 = _T_378 ? _GEN_144 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 697:9:@5881.20]
  assign _GEN_150 = _T_378 ? _GEN_145 : blockCounter; // @[pageswappergcm.scala 697:9:@5881.20]
  assign _GEN_151 = _T_823 ? 1'h0 : tagUp; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_152 = _T_823 ? _GEN_130 : _GEN_149; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_153 = _T_823 ? tagState : _GEN_146; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_154 = _T_823 ? cleanupStateNext : _GEN_147; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_155 = _T_823 ? _GEN_101 : _GEN_148; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_156 = _T_823 ? blockCounter : _GEN_150; // @[pageswappergcm.scala 684:9:@5870.18]
  assign _GEN_161 = _T_462 ? _GEN_124 : _GEN_106; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_162 = _T_462 ? _GEN_125 : _GEN_107; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_163 = _T_462 ? _GEN_126 : _GEN_108; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_164 = _T_462 ? _GEN_127 : _GEN_109; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_165 = _T_462 ? _GEN_128 : _GEN_151; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_166 = _T_462 ? {{7'd0}, _GEN_129} : _GEN_152; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_167 = _T_462 ? tagState : _GEN_153; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_168 = _T_462 ? cleanupStateNext : _GEN_154; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_169 = _T_462 ? _GEN_101 : _GEN_155; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_170 = _T_462 ? blockCounter : _GEN_156; // @[pageswappergcm.scala 629:9:@5844.16]
  assign _GEN_171 = _T_283 ? {{7'd0}, _T_798} : _GEN_166; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_172 = _T_283 ? _GEN_119 : _GEN_170; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_173 = _T_283 ? 2'h2 : _GEN_167; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_178 = _T_283 ? _GEN_106 : _GEN_161; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_179 = _T_283 ? _GEN_107 : _GEN_162; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_180 = _T_283 ? _GEN_108 : _GEN_163; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_181 = _T_283 ? _GEN_109 : _GEN_164; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_182 = _T_283 ? tagUp : _GEN_165; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_183 = _T_283 ? cleanupStateNext : _GEN_168; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_184 = _T_283 ? _GEN_101 : _GEN_169; // @[pageswappergcm.scala 602:9:@5820.14]
  assign _GEN_185 = cond1 ? _GEN_115 : _GEN_103; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_186 = cond1 ? _GEN_116 : _GEN_183; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_187 = cond1 ? {{7'd0}, _GEN_110} : _GEN_171; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_188 = cond1 ? blockCounter : _GEN_172; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_189 = cond1 ? tagState : _GEN_173; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_194 = cond1 ? _GEN_106 : _GEN_178; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_195 = cond1 ? _GEN_107 : _GEN_179; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_196 = cond1 ? _GEN_108 : _GEN_180; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_197 = cond1 ? _GEN_109 : _GEN_181; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_198 = cond1 ? tagUp : _GEN_182; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_199 = cond1 ? _GEN_101 : _GEN_184; // @[pageswappergcm.scala 591:9:@5811.12]
  assign _GEN_200 = _T_290 ? {{4'd0}, _T_787} : _GEN_187; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_201 = _T_290 ? _GEN_103 : _GEN_185; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_202 = _T_290 ? cleanupStateNext : _GEN_186; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_203 = _T_290 ? blockCounter : _GEN_188; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_204 = _T_290 ? tagState : _GEN_189; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_209 = _T_290 ? _GEN_106 : _GEN_194; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_210 = _T_290 ? _GEN_107 : _GEN_195; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_211 = _T_290 ? _GEN_108 : _GEN_196; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_212 = _T_290 ? _GEN_109 : _GEN_197; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_213 = _T_290 ? tagUp : _GEN_198; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_214 = _T_290 ? _GEN_101 : _GEN_199; // @[pageswappergcm.scala 586:9:@5803.10]
  assign _GEN_215 = _T_629 ? 32'h20 : _GEN_103; // @[pageswappergcm.scala 736:13:@5924.14]
  assign _GEN_216 = _T_629 ? 2'h0 : cleanupStateNext; // @[pageswappergcm.scala 736:13:@5924.14]
  assign _T_868 = 39'h1 << 3'h5; // @[pageswappergcm.scala 749:53:@5938.20]
  assign _T_869 = ~ _T_868; // @[pageswappergcm.scala 749:42:@5939.20]
  assign _T_870 = _GEN_443 & _T_869; // @[pageswappergcm.scala 749:40:@5940.20]
  assign _GEN_217 = pindataReady ? _T_870 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 748:13:@5937.18]
  assign _GEN_218 = pindataReady ? 3'h2 : _T_774; // @[pageswappergcm.scala 748:13:@5937.18]
  assign _GEN_219 = aesm_io_newR ? _T_810 : _GEN_111; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _GEN_220 = aesm_io_newR ? _T_811 : _GEN_112; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _GEN_221 = aesm_io_newR ? _T_812 : _GEN_113; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _GEN_222 = aesm_io_newR ? _T_813 : _GEN_114; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _GEN_223 = aesm_io_newR ? 3'h3 : _T_774; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _GEN_225 = aesm_io_newR ? _T_803 : blockCounter; // @[pageswappergcm.scala 755:13:@5948.20]
  assign _T_890 = blockCounter - 32'h1; // @[pageswappergcm.scala 776:33:@5973.22]
  assign _T_891 = $unsigned(_T_890); // @[pageswappergcm.scala 776:33:@5974.22]
  assign _T_892 = _T_891[31:0]; // @[pageswappergcm.scala 776:33:@5975.22]
  assign _T_894 = _T_892 == 32'h0; // @[pageswappergcm.scala 776:39:@5976.22]
  assign _T_901 = _T_892 < ConfReg_2; // @[pageswappergcm.scala 792:45:@5987.28]
  assign _GEN_226 = _T_901 ? 3'h1 : 3'h5; // @[pageswappergcm.scala 793:21:@5988.28]
  assign _GEN_227 = io_memio_ready ? _GEN_226 : _T_774; // @[pageswappergcm.scala 790:19:@5983.26]
  assign _GEN_229 = _T_627 ? _GEN_227 : _GEN_226; // @[pageswappergcm.scala 782:17:@5982.24]
  assign _GEN_230 = _T_894 ? 3'h2 : _GEN_229; // @[pageswappergcm.scala 777:15:@5977.22]
  assign _T_926 = _T_844 & _T_869; // @[pageswappergcm.scala 829:59:@6034.30]
  assign _T_929 = sessionIv == tag; // @[pageswappergcm.scala 842:30:@6040.30]
  assign _T_932 = ConfReg_4 & 32'h1; // @[pageswappergcm.scala 844:42:@6043.32]
  assign _T_934 = ConfReg_4 | 32'h2; // @[pageswappergcm.scala 847:42:@6047.32]
  assign _GEN_231 = _T_929 ? _T_932 : _T_934; // @[pageswappergcm.scala 843:15:@6041.30]
  assign _GEN_233 = _T_311 ? _T_926 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 826:12:@6027.28]
  assign _GEN_234 = _T_311 ? 3'h6 : _T_774; // @[pageswappergcm.scala 826:12:@6027.28]
  assign _GEN_238 = _T_311 ? _GEN_231 : _T_700; // @[pageswappergcm.scala 826:12:@6027.28]
  assign _GEN_242 = _T_835 ? {{7'd0}, _GEN_110} : _GEN_233; // @[pageswappergcm.scala 822:12:@6021.26]
  assign _GEN_243 = _T_835 ? _T_774 : _GEN_234; // @[pageswappergcm.scala 822:12:@6021.26]
  assign _GEN_245 = _T_835 ? _T_700 : _GEN_238; // @[pageswappergcm.scala 822:12:@6021.26]
  assign _GEN_249 = _T_263 ? {{7'd0}, _GEN_110} : _GEN_242; // @[pageswappergcm.scala 817:12:@6016.24]
  assign _GEN_250 = _T_263 ? _T_774 : _GEN_243; // @[pageswappergcm.scala 817:12:@6016.24]
  assign _GEN_252 = _T_263 ? _T_700 : _GEN_245; // @[pageswappergcm.scala 817:12:@6016.24]
  assign _GEN_256 = _T_378 ? _GEN_249 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 810:11:@6013.22]
  assign _GEN_257 = _T_378 ? _GEN_250 : _T_774; // @[pageswappergcm.scala 810:11:@6013.22]
  assign _GEN_259 = _T_378 ? _GEN_252 : _T_700; // @[pageswappergcm.scala 810:11:@6013.22]
  assign _GEN_260 = _T_436 ? {{4'd0}, _T_787} : _GEN_256; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_261 = _T_436 ? _GEN_230 : _GEN_257; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_262 = _T_436 ? 2'h2 : _GEN_146; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_263 = _T_436 ? cleanupStateNext : _GEN_147; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_264 = _T_436 ? _GEN_101 : _GEN_148; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_265 = _T_436 ? blockCounter : _GEN_150; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_266 = _T_436 ? _T_700 : _GEN_259; // @[pageswappergcm.scala 774:11:@5968.20]
  assign _GEN_267 = _T_462 ? _GEN_219 : _GEN_111; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_268 = _T_462 ? _GEN_220 : _GEN_112; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_269 = _T_462 ? _GEN_221 : _GEN_113; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_270 = _T_462 ? _GEN_222 : _GEN_114; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_271 = _T_462 ? _GEN_223 : _GEN_261; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_272 = _T_462 ? {{7'd0}, _GEN_129} : _GEN_260; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_273 = _T_462 ? _GEN_225 : _GEN_265; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_274 = _T_462 ? tagState : _GEN_262; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_275 = _T_462 ? cleanupStateNext : _GEN_263; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_276 = _T_462 ? _GEN_101 : _GEN_264; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_277 = _T_462 ? _T_700 : _GEN_266; // @[pageswappergcm.scala 753:11:@5947.18]
  assign _GEN_278 = _T_283 ? _GEN_217 : _GEN_272; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_279 = _T_283 ? _GEN_218 : _GEN_271; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_280 = _T_283 ? _GEN_111 : _GEN_267; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_281 = _T_283 ? _GEN_112 : _GEN_268; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_282 = _T_283 ? _GEN_113 : _GEN_269; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_283 = _T_283 ? _GEN_114 : _GEN_270; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_284 = _T_283 ? blockCounter : _GEN_273; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_285 = _T_283 ? tagState : _GEN_274; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_286 = _T_283 ? cleanupStateNext : _GEN_275; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_287 = _T_283 ? _GEN_101 : _GEN_276; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_288 = _T_283 ? _T_700 : _GEN_277; // @[pageswappergcm.scala 746:11:@5936.16]
  assign _GEN_289 = cond1 ? 3'h1 : _GEN_279; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_290 = cond1 ? {{7'd0}, _GEN_110} : _GEN_278; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_291 = cond1 ? _GEN_111 : _GEN_280; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_292 = cond1 ? _GEN_112 : _GEN_281; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_293 = cond1 ? _GEN_113 : _GEN_282; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_294 = cond1 ? _GEN_114 : _GEN_283; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_295 = cond1 ? blockCounter : _GEN_284; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_296 = cond1 ? tagState : _GEN_285; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_297 = cond1 ? cleanupStateNext : _GEN_286; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_298 = cond1 ? _GEN_101 : _GEN_287; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_299 = cond1 ? _T_700 : _GEN_288; // @[pageswappergcm.scala 743:11:@5931.14]
  assign _GEN_300 = _T_290 ? 3'h0 : _GEN_289; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_301 = _T_290 ? {{4'd0}, _T_787} : _GEN_290; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_302 = _T_290 ? _GEN_215 : _GEN_103; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_303 = _T_290 ? _GEN_216 : _GEN_297; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_304 = _T_290 ? _GEN_111 : _GEN_291; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_305 = _T_290 ? _GEN_112 : _GEN_292; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_306 = _T_290 ? _GEN_113 : _GEN_293; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_307 = _T_290 ? _GEN_114 : _GEN_294; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_308 = _T_290 ? blockCounter : _GEN_295; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_309 = _T_290 ? tagState : _GEN_296; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_310 = _T_290 ? _GEN_101 : _GEN_298; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_311 = _T_290 ? _T_700 : _GEN_299; // @[pageswappergcm.scala 731:11:@5917.12]
  assign _GEN_312 = _T_630 ? _GEN_300 : _T_774; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_313 = _T_630 ? _GEN_301 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_314 = _T_630 ? _GEN_302 : _GEN_103; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_315 = _T_630 ? _GEN_303 : cleanupStateNext; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_316 = _T_630 ? _GEN_304 : _GEN_111; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_317 = _T_630 ? _GEN_305 : _GEN_112; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_318 = _T_630 ? _GEN_306 : _GEN_113; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_319 = _T_630 ? _GEN_307 : _GEN_114; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_320 = _T_630 ? _GEN_308 : blockCounter; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_321 = _T_630 ? _GEN_309 : tagState; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_322 = _T_630 ? _GEN_310 : _GEN_101; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_323 = _T_630 ? _GEN_311 : _T_700; // @[pageswappergcm.scala 729:7:@5915.10]
  assign _GEN_324 = _T_222 ? _GEN_200 : _GEN_313; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_325 = _T_222 ? _GEN_201 : _GEN_314; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_326 = _T_222 ? _GEN_202 : _GEN_315; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_327 = _T_222 ? _GEN_203 : _GEN_320; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_328 = _T_222 ? _GEN_204 : _GEN_321; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_333 = _T_222 ? _GEN_209 : _GEN_106; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_334 = _T_222 ? _GEN_210 : _GEN_107; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_335 = _T_222 ? _GEN_211 : _GEN_108; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_336 = _T_222 ? _GEN_212 : _GEN_109; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_337 = _T_222 ? _GEN_213 : tagUp; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_338 = _T_222 ? _GEN_214 : _GEN_322; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_339 = _T_222 ? _T_774 : _GEN_312; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_340 = _T_222 ? _GEN_111 : _GEN_316; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_341 = _T_222 ? _GEN_112 : _GEN_317; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_342 = _T_222 ? _GEN_113 : _GEN_318; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_343 = _T_222 ? _GEN_114 : _GEN_319; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_344 = _T_222 ? _T_700 : _GEN_323; // @[pageswappergcm.scala 583:7:@5801.8]
  assign _GEN_345 = start ? _GEN_324 : {{7'd0}, _GEN_110}; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_346 = start ? _GEN_325 : _GEN_103; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_347 = start ? _GEN_326 : cleanupStateNext; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_348 = start ? _GEN_327 : blockCounter; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_349 = start ? _GEN_328 : tagState; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_354 = start ? _GEN_333 : _GEN_106; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_355 = start ? _GEN_334 : _GEN_107; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_356 = start ? _GEN_335 : _GEN_108; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_357 = start ? _GEN_336 : _GEN_109; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_358 = start ? _GEN_337 : tagUp; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_359 = start ? _GEN_338 : _GEN_101; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_360 = start ? _GEN_339 : _T_774; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_361 = start ? _GEN_340 : _GEN_111; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_362 = start ? _GEN_341 : _GEN_112; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_363 = start ? _GEN_342 : _GEN_113; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_364 = start ? _GEN_343 : _GEN_114; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _GEN_365 = start ? _GEN_344 : _T_700; // @[pageswappergcm.scala 580:5:@5797.6]
  assign _T_937 = initState == 3'h0; // @[pageswappergcm.scala 862:20:@6060.6]
  assign _T_938 = initState == 3'h1; // @[pageswappergcm.scala 865:26:@6065.8]
  assign _GEN_366 = rndgenm_io_done ? rndgenm_io_out : nonce; // @[pageswappergcm.scala 868:11:@6067.10]
  assign _GEN_367 = rndgenm_io_done ? 3'h2 : initStateNext; // @[pageswappergcm.scala 868:11:@6067.10]
  assign _T_939 = initState == 3'h2; // @[pageswappergcm.scala 872:26:@6073.10]
  assign _GEN_368 = rndgenm_io_done ? {{64'd0}, rndgenm_io_out} : sessionKey; // @[pageswappergcm.scala 875:11:@6075.12]
  assign _GEN_369 = rndgenm_io_done ? 3'h3 : initStateNext; // @[pageswappergcm.scala 875:11:@6075.12]
  assign _T_940 = initState == 3'h3; // @[pageswappergcm.scala 879:26:@6081.12]
  assign _GEN_450 = {{127'd0}, rndgenm_io_out}; // @[pageswappergcm.scala 883:51:@6084.16]
  assign _T_942 = _GEN_450 << 7'h40; // @[pageswappergcm.scala 883:51:@6084.16]
  assign _GEN_451 = {{63'd0}, sessionKey}; // @[pageswappergcm.scala 883:34:@6085.16]
  assign _T_943 = _GEN_451 | _T_942; // @[pageswappergcm.scala 883:34:@6085.16]
  assign _GEN_370 = rndgenm_io_done ? _T_943 : {{63'd0}, sessionKey}; // @[pageswappergcm.scala 882:11:@6083.14]
  assign _GEN_371 = rndgenm_io_done ? 3'h4 : initStateNext; // @[pageswappergcm.scala 882:11:@6083.14]
  assign _GEN_372 = rndgenm_io_done ? 3'h5 : initStateNext; // @[pageswappergcm.scala 890:9:@6093.16]
  assign _T_948 = 2'h1 << 1'h1; // @[pageswappergcm.scala 903:46:@6102.20]
  assign _GEN_452 = {{30'd0}, _T_948}; // @[pageswappergcm.scala 903:40:@6103.20]
  assign _T_949 = ConfReg_9 | _GEN_452; // @[pageswappergcm.scala 903:40:@6103.20]
  assign _GEN_373 = aesm_io_newR ? aesm_io_out : h; // @[pageswappergcm.scala 896:11:@6100.18]
  assign _GEN_374 = aesm_io_newR ? _T_949 : _GEN_110; // @[pageswappergcm.scala 896:11:@6100.18]
  assign _GEN_375 = aesm_io_newR ? 3'h6 : initStateNext; // @[pageswappergcm.scala 896:11:@6100.18]
  assign _GEN_376 = _T_522 ? _GEN_373 : h; // @[pageswappergcm.scala 894:6:@6099.16]
  assign _GEN_377 = _T_522 ? _GEN_374 : _GEN_110; // @[pageswappergcm.scala 894:6:@6099.16]
  assign _GEN_378 = _T_522 ? _GEN_375 : initStateNext; // @[pageswappergcm.scala 894:6:@6099.16]
  assign _GEN_379 = _T_274 ? _GEN_372 : _GEN_378; // @[pageswappergcm.scala 888:6:@6092.14]
  assign _GEN_380 = _T_274 ? h : _GEN_376; // @[pageswappergcm.scala 888:6:@6092.14]
  assign _GEN_381 = _T_274 ? _GEN_110 : _GEN_377; // @[pageswappergcm.scala 888:6:@6092.14]
  assign _GEN_382 = _T_940 ? _GEN_370 : {{63'd0}, sessionKey}; // @[pageswappergcm.scala 880:5:@6082.12]
  assign _GEN_383 = _T_940 ? _GEN_371 : _GEN_379; // @[pageswappergcm.scala 880:5:@6082.12]
  assign _GEN_384 = _T_940 ? h : _GEN_380; // @[pageswappergcm.scala 880:5:@6082.12]
  assign _GEN_385 = _T_940 ? _GEN_110 : _GEN_381; // @[pageswappergcm.scala 880:5:@6082.12]
  assign _GEN_386 = _T_939 ? {{63'd0}, _GEN_368} : _GEN_382; // @[pageswappergcm.scala 873:5:@6074.10]
  assign _GEN_387 = _T_939 ? _GEN_369 : _GEN_383; // @[pageswappergcm.scala 873:5:@6074.10]
  assign _GEN_388 = _T_939 ? h : _GEN_384; // @[pageswappergcm.scala 873:5:@6074.10]
  assign _GEN_389 = _T_939 ? _GEN_110 : _GEN_385; // @[pageswappergcm.scala 873:5:@6074.10]
  assign _GEN_390 = _T_938 ? _GEN_366 : nonce; // @[pageswappergcm.scala 866:5:@6066.8]
  assign _GEN_391 = _T_938 ? _GEN_367 : _GEN_387; // @[pageswappergcm.scala 866:5:@6066.8]
  assign _GEN_392 = _T_938 ? {{63'd0}, sessionKey} : _GEN_386; // @[pageswappergcm.scala 866:5:@6066.8]
  assign _GEN_393 = _T_938 ? h : _GEN_388; // @[pageswappergcm.scala 866:5:@6066.8]
  assign _GEN_394 = _T_938 ? _GEN_110 : _GEN_389; // @[pageswappergcm.scala 866:5:@6066.8]
  assign _GEN_395 = _T_937 ? 3'h1 : _GEN_391; // @[pageswappergcm.scala 863:5:@6061.6]
  assign _GEN_396 = _T_937 ? nonce : _GEN_390; // @[pageswappergcm.scala 863:5:@6061.6]
  assign _GEN_397 = _T_937 ? {{63'd0}, sessionKey} : _GEN_392; // @[pageswappergcm.scala 863:5:@6061.6]
  assign _GEN_398 = _T_937 ? h : _GEN_393; // @[pageswappergcm.scala 863:5:@6061.6]
  assign _GEN_399 = _T_937 ? _GEN_110 : _GEN_394; // @[pageswappergcm.scala 863:5:@6061.6]
  assign _GEN_400 = moduleReady ? _GEN_345 : {{7'd0}, _GEN_399}; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_401 = moduleReady ? _GEN_346 : _GEN_103; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_402 = moduleReady ? _GEN_347 : cleanupStateNext; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_403 = moduleReady ? _GEN_348 : blockCounter; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_404 = moduleReady ? _GEN_349 : tagState; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_409 = moduleReady ? _GEN_354 : _GEN_106; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_410 = moduleReady ? _GEN_355 : _GEN_107; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_411 = moduleReady ? _GEN_356 : _GEN_108; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_412 = moduleReady ? _GEN_357 : _GEN_109; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_413 = moduleReady ? _GEN_358 : tagUp; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_414 = moduleReady ? _GEN_359 : _GEN_101; // @[pageswappergcm.scala 576:3:@5795.4]
  assign poStateNext = moduleReady ? _GEN_360 : _T_774; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_416 = moduleReady ? _GEN_361 : _GEN_111; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_417 = moduleReady ? _GEN_362 : _GEN_112; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_418 = moduleReady ? _GEN_363 : _GEN_113; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_419 = moduleReady ? _GEN_364 : _GEN_114; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_420 = moduleReady ? _GEN_365 : _T_700; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_421 = moduleReady ? initStateNext : _GEN_395; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_422 = moduleReady ? nonce : _GEN_396; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_423 = moduleReady ? {{63'd0}, sessionKey} : _GEN_397; // @[pageswappergcm.scala 576:3:@5795.4]
  assign _GEN_424 = moduleReady ? h : _GEN_398; // @[pageswappergcm.scala 576:3:@5795.4]
  assign io_mainMemio_rdata = _T_608;
  assign io_mainMemio_ready = _T_620;
  assign io_socMemio_addr = io_mainMemio_addr;
  assign io_socMemio_wdata = io_mainMemio_wdata;
  assign io_socMemio_we = _T_598;
  assign io_socMemio_en = _T_603;
  assign io_memio_addr = addr[10:0];
  assign io_memio_wdata = _T_748;
  assign io_memio_we = _T_300;
  assign io_memio_en = mmenvalid;
  assign io_err = _T_497;
  assign io_currOutReady = _T_495;
  assign io_finished = _T_498;
  assign rndgenm_clock = clock;
  assign rndgenm_reset = reset;
  assign rndgenm_io_en = _T_270;
  assign cntrm_clock = clock;
  assign cntrm_io_get = newC;
  assign cntrm_io_reset = _T_275;
  assign cntrm_io_init = _T_281;
  assign vfm_clock = clock;
  assign vfm_reset = reset;
  assign vfm_io_wdata = _T_428[256:0];
  assign vfm_io_addr = _T_395[4:0];
  assign vfm_io_cmd = _T_376;
  assign aesm_clock = clock;
  assign aesm_reset = reset;
  assign aesm_io_intVect = _T_528;
  assign aesm_io_data = _T_556;
  assign aesm_io_en = encry;
  assign aesm_io_key = sessionKey;
  assign gmultm_io_x = h;
  assign gmultm_io_y = _T_249;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{$random}};
  h = _RAND_0[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {4{$random}};
  tag = _RAND_1[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {4{$random}};
  IVTag = _RAND_2[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {2{$random}};
  nonce = _RAND_3[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {4{$random}};
  curriv = _RAND_4[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {4{$random}};
  sessionIv = _RAND_5[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {4{$random}};
  sessionKey = _RAND_6[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  blockCounter = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {4{$random}};
  currBlockBuff = _RAND_8[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  ConfReg_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  ConfReg_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  ConfReg_2 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  ConfReg_3 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  ConfReg_4 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  ConfReg_5 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  ConfReg_6 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  ConfReg_7 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  ConfReg_8 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  ConfReg_9 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  ConfReg_10 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  ConfReg_11 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  ConfReg_12 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  ConfReg_13 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  initState = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  initStateNext = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  poState = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  cleanupState = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  cleanupStateNext = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  tagState = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  tagUp = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  encry = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      h <= 128'h0;
    end else begin
      if (!(moduleReady)) begin
        if (!(_T_937)) begin
          if (!(_T_938)) begin
            if (!(_T_939)) begin
              if (!(_T_940)) begin
                if (!(_T_274)) begin
                  if (_T_522) begin
                    if (aesm_io_newR) begin
                      h <= aesm_io_out;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tag <= 128'h0;
    end else begin
      if (_T_246) begin
        if (_T_260) begin
          tag <= gmultm_io_out;
        end
      end else begin
        if (_T_244) begin
          if (_T_263) begin
            tag <= gmultm_io_out;
          end else begin
            tag <= _T_264;
          end
        end
      end
    end
    if (reset) begin
      IVTag <= 128'h0;
    end else begin
      if (_T_251) begin
        IVTag <= 128'h0;
      end else begin
        if (_T_253) begin
          if (aesDone) begin
            if (_T_222) begin
              IVTag <= aesdecInput;
            end else begin
              IVTag <= _T_225;
            end
          end else begin
            IVTag <= 128'h0;
          end
        end
      end
    end
    if (reset) begin
      nonce <= 64'h0;
    end else begin
      if (!(moduleReady)) begin
        if (!(_T_937)) begin
          if (_T_938) begin
            if (rndgenm_io_done) begin
              nonce <= rndgenm_io_out;
            end
          end
        end
      end
    end
    if (reset) begin
      curriv <= 128'h0;
    end else begin
      curriv <= xcv[127:0];
    end
    if (reset) begin
      sessionIv <= 128'h0;
    end else begin
      sessionIv <= _T_474[127:0];
    end
    if (reset) begin
      sessionKey <= 128'h0;
    end else begin
      sessionKey <= _GEN_423[127:0];
    end
    if (reset) begin
      blockCounter <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (!(_T_290)) begin
              if (!(cond1)) begin
                if (_T_283) begin
                  if (_T_219) begin
                    if (io_memio_ready) begin
                      blockCounter <= _T_803;
                    end
                  end else begin
                    if (_T_221) begin
                      blockCounter <= _T_803;
                    end
                  end
                end else begin
                  if (!(_T_462)) begin
                    if (!(_T_823)) begin
                      if (_T_378) begin
                        if (!(_T_263)) begin
                          if (!(_T_835)) begin
                            if (_T_311) begin
                              blockCounter <= 32'h0;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (!(_T_290)) begin
                if (!(cond1)) begin
                  if (!(_T_283)) begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        blockCounter <= _T_803;
                      end
                    end else begin
                      if (!(_T_436)) begin
                        if (_T_378) begin
                          if (!(_T_263)) begin
                            if (!(_T_835)) begin
                              if (_T_311) begin
                                blockCounter <= 32'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      currBlockBuff <= 128'h0;
    end else begin
      if (_T_304) begin
        if (_T_253) begin
          currBlockBuff <= 128'h0;
        end else begin
          if (_T_283) begin
            currBlockBuff <= io_memio_rdata;
          end
        end
      end else begin
        if (_T_302) begin
          if (_T_253) begin
            currBlockBuff <= 128'h0;
          end else begin
            currBlockBuff <= vfm_io_rdata;
          end
        end else begin
          if (_T_300) begin
            currBlockBuff <= aesdecInput;
          end else begin
            if (_T_298) begin
              currBlockBuff <= aesdecInput;
            end
          end
        end
      end
    end
    if (reset) begin
      ConfReg_0 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h0 == confaddr) begin
                        ConfReg_0 <= _T_656;
                      end
                    end else begin
                      if (4'h0 == confaddr) begin
                        ConfReg_0 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h0 == confaddr) begin
                          ConfReg_0 <= _T_656;
                        end
                      end else begin
                        if (4'h0 == confaddr) begin
                          ConfReg_0 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_283) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h0 == confaddr) begin
                            ConfReg_0 <= _T_656;
                          end
                        end else begin
                          if (4'h0 == confaddr) begin
                            ConfReg_0 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_462) begin
                    if (_T_611) begin
                      if (_T_642) begin
                        if (io_mainMemio_we) begin
                          if (_T_647) begin
                            if (4'h0 == confaddr) begin
                              ConfReg_0 <= _T_656;
                            end
                          end else begin
                            if (4'h0 == confaddr) begin
                              ConfReg_0 <= _T_644;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_823) begin
                      ConfReg_0 <= _GEN_101;
                    end else begin
                      if (_T_378) begin
                        if (_T_263) begin
                          ConfReg_0 <= _GEN_101;
                        end else begin
                          if (_T_835) begin
                            ConfReg_0 <= _GEN_101;
                          end else begin
                            if (_T_311) begin
                              ConfReg_0 <= _T_840;
                            end else begin
                              ConfReg_0 <= _GEN_101;
                            end
                          end
                        end
                      end else begin
                        ConfReg_0 <= _GEN_101;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                ConfReg_0 <= _GEN_101;
              end else begin
                if (cond1) begin
                  ConfReg_0 <= _GEN_101;
                end else begin
                  if (_T_283) begin
                    ConfReg_0 <= _GEN_101;
                  end else begin
                    if (_T_462) begin
                      ConfReg_0 <= _GEN_101;
                    end else begin
                      if (_T_436) begin
                        ConfReg_0 <= _GEN_101;
                      end else begin
                        if (_T_378) begin
                          if (_T_263) begin
                            ConfReg_0 <= _GEN_101;
                          end else begin
                            if (_T_835) begin
                              ConfReg_0 <= _GEN_101;
                            end else begin
                              if (_T_311) begin
                                ConfReg_0 <= _T_840;
                              end else begin
                                ConfReg_0 <= _GEN_101;
                              end
                            end
                          end
                        end else begin
                          ConfReg_0 <= _GEN_101;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              ConfReg_0 <= _GEN_101;
            end
          end
        end else begin
          ConfReg_0 <= _GEN_101;
        end
      end else begin
        ConfReg_0 <= _GEN_101;
      end
    end
    if (reset) begin
      ConfReg_1 <= 32'h0;
    end else begin
      if (_T_611) begin
        if (_T_642) begin
          if (io_mainMemio_we) begin
            if (_T_647) begin
              if (4'h1 == confaddr) begin
                ConfReg_1 <= _T_656;
              end
            end else begin
              if (4'h1 == confaddr) begin
                ConfReg_1 <= _T_644;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      ConfReg_2 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h2 == confaddr) begin
                        ConfReg_2 <= _T_656;
                      end
                    end else begin
                      if (4'h2 == confaddr) begin
                        ConfReg_2 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_221) begin
                  ConfReg_2 <= 32'h20;
                end else begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h2 == confaddr) begin
                            ConfReg_2 <= _T_656;
                          end
                        end else begin
                          if (4'h2 == confaddr) begin
                            ConfReg_2 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h2 == confaddr) begin
                          ConfReg_2 <= _T_656;
                        end
                      end else begin
                        if (4'h2 == confaddr) begin
                          ConfReg_2 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_629) begin
                  ConfReg_2 <= 32'h20;
                end else begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h2 == confaddr) begin
                            ConfReg_2 <= _T_656;
                          end
                        end else begin
                          if (4'h2 == confaddr) begin
                            ConfReg_2 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end
              end else begin
                ConfReg_2 <= _GEN_103;
              end
            end else begin
              ConfReg_2 <= _GEN_103;
            end
          end
        end else begin
          ConfReg_2 <= _GEN_103;
        end
      end else begin
        ConfReg_2 <= _GEN_103;
      end
    end
    if (reset) begin
      ConfReg_3 <= 32'h0;
    end else begin
      ConfReg_3 <= _T_689[31:0];
    end
    if (reset) begin
      ConfReg_4 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (start) begin
              if (_T_304) begin
                if (_T_694) begin
                  ConfReg_4 <= _T_696;
                end
              end else begin
                ConfReg_4 <= 32'h0;
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (start) begin
                  if (_T_304) begin
                    if (_T_694) begin
                      ConfReg_4 <= _T_696;
                    end
                  end else begin
                    ConfReg_4 <= 32'h0;
                  end
                end
              end else begin
                if (cond1) begin
                  if (start) begin
                    if (_T_304) begin
                      if (_T_694) begin
                        ConfReg_4 <= _T_696;
                      end
                    end else begin
                      ConfReg_4 <= 32'h0;
                    end
                  end
                end else begin
                  if (_T_283) begin
                    if (start) begin
                      if (_T_304) begin
                        if (_T_694) begin
                          ConfReg_4 <= _T_696;
                        end
                      end else begin
                        ConfReg_4 <= 32'h0;
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      ConfReg_4 <= _T_700;
                    end else begin
                      if (_T_436) begin
                        ConfReg_4 <= _T_700;
                      end else begin
                        if (_T_378) begin
                          if (_T_263) begin
                            ConfReg_4 <= _T_700;
                          end else begin
                            if (_T_835) begin
                              ConfReg_4 <= _T_700;
                            end else begin
                              if (_T_311) begin
                                if (_T_929) begin
                                  ConfReg_4 <= _T_932;
                                end else begin
                                  ConfReg_4 <= _T_934;
                                end
                              end else begin
                                ConfReg_4 <= _T_700;
                              end
                            end
                          end
                        end else begin
                          ConfReg_4 <= _T_700;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              ConfReg_4 <= _T_700;
            end
          end
        end else begin
          ConfReg_4 <= _T_700;
        end
      end else begin
        ConfReg_4 <= _T_700;
      end
    end
    if (reset) begin
      ConfReg_5 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h5 == confaddr) begin
                        ConfReg_5 <= _T_656;
                      end
                    end else begin
                      if (4'h5 == confaddr) begin
                        ConfReg_5 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h5 == confaddr) begin
                          ConfReg_5 <= _T_656;
                        end
                      end else begin
                        if (4'h5 == confaddr) begin
                          ConfReg_5 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_283) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h5 == confaddr) begin
                            ConfReg_5 <= _T_656;
                          end
                        end else begin
                          if (4'h5 == confaddr) begin
                            ConfReg_5 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_462) begin
                    if (aesm_io_newR) begin
                      ConfReg_5 <= _T_810;
                    end else begin
                      if (_T_611) begin
                        if (_T_642) begin
                          if (io_mainMemio_we) begin
                            if (_T_647) begin
                              if (4'h5 == confaddr) begin
                                ConfReg_5 <= _T_656;
                              end
                            end else begin
                              if (4'h5 == confaddr) begin
                                ConfReg_5 <= _T_644;
                              end
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    ConfReg_5 <= _GEN_106;
                  end
                end
              end
            end
          end else begin
            ConfReg_5 <= _GEN_106;
          end
        end else begin
          ConfReg_5 <= _GEN_106;
        end
      end else begin
        ConfReg_5 <= _GEN_106;
      end
    end
    if (reset) begin
      ConfReg_6 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h6 == confaddr) begin
                        ConfReg_6 <= _T_656;
                      end
                    end else begin
                      if (4'h6 == confaddr) begin
                        ConfReg_6 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h6 == confaddr) begin
                          ConfReg_6 <= _T_656;
                        end
                      end else begin
                        if (4'h6 == confaddr) begin
                          ConfReg_6 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_283) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h6 == confaddr) begin
                            ConfReg_6 <= _T_656;
                          end
                        end else begin
                          if (4'h6 == confaddr) begin
                            ConfReg_6 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_462) begin
                    if (aesm_io_newR) begin
                      ConfReg_6 <= _T_811;
                    end else begin
                      if (_T_611) begin
                        if (_T_642) begin
                          if (io_mainMemio_we) begin
                            if (_T_647) begin
                              if (4'h6 == confaddr) begin
                                ConfReg_6 <= _T_656;
                              end
                            end else begin
                              if (4'h6 == confaddr) begin
                                ConfReg_6 <= _T_644;
                              end
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    ConfReg_6 <= _GEN_107;
                  end
                end
              end
            end
          end else begin
            ConfReg_6 <= _GEN_107;
          end
        end else begin
          ConfReg_6 <= _GEN_107;
        end
      end else begin
        ConfReg_6 <= _GEN_107;
      end
    end
    if (reset) begin
      ConfReg_7 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h7 == confaddr) begin
                        ConfReg_7 <= _T_656;
                      end
                    end else begin
                      if (4'h7 == confaddr) begin
                        ConfReg_7 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h7 == confaddr) begin
                          ConfReg_7 <= _T_656;
                        end
                      end else begin
                        if (4'h7 == confaddr) begin
                          ConfReg_7 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_283) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h7 == confaddr) begin
                            ConfReg_7 <= _T_656;
                          end
                        end else begin
                          if (4'h7 == confaddr) begin
                            ConfReg_7 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_462) begin
                    if (aesm_io_newR) begin
                      ConfReg_7 <= _T_812;
                    end else begin
                      if (_T_611) begin
                        if (_T_642) begin
                          if (io_mainMemio_we) begin
                            if (_T_647) begin
                              if (4'h7 == confaddr) begin
                                ConfReg_7 <= _T_656;
                              end
                            end else begin
                              if (4'h7 == confaddr) begin
                                ConfReg_7 <= _T_644;
                              end
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    ConfReg_7 <= _GEN_108;
                  end
                end
              end
            end
          end else begin
            ConfReg_7 <= _GEN_108;
          end
        end else begin
          ConfReg_7 <= _GEN_108;
        end
      end else begin
        ConfReg_7 <= _GEN_108;
      end
    end
    if (reset) begin
      ConfReg_8 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_290) begin
              if (_T_611) begin
                if (_T_642) begin
                  if (io_mainMemio_we) begin
                    if (_T_647) begin
                      if (4'h8 == confaddr) begin
                        ConfReg_8 <= _T_656;
                      end
                    end else begin
                      if (4'h8 == confaddr) begin
                        ConfReg_8 <= _T_644;
                      end
                    end
                  end
                end
              end
            end else begin
              if (cond1) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'h8 == confaddr) begin
                          ConfReg_8 <= _T_656;
                        end
                      end else begin
                        if (4'h8 == confaddr) begin
                          ConfReg_8 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_283) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'h8 == confaddr) begin
                            ConfReg_8 <= _T_656;
                          end
                        end else begin
                          if (4'h8 == confaddr) begin
                            ConfReg_8 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_462) begin
                    if (aesm_io_newR) begin
                      ConfReg_8 <= _T_813;
                    end else begin
                      if (_T_611) begin
                        if (_T_642) begin
                          if (io_mainMemio_we) begin
                            if (_T_647) begin
                              if (4'h8 == confaddr) begin
                                ConfReg_8 <= _T_656;
                              end
                            end else begin
                              if (4'h8 == confaddr) begin
                                ConfReg_8 <= _T_644;
                              end
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    ConfReg_8 <= _GEN_109;
                  end
                end
              end
            end
          end else begin
            ConfReg_8 <= _GEN_109;
          end
        end else begin
          ConfReg_8 <= _GEN_109;
        end
      end else begin
        ConfReg_8 <= _GEN_109;
      end
    end
    if (reset) begin
      ConfReg_9 <= 32'h0;
    end else begin
      ConfReg_9 <= _GEN_400[31:0];
    end
    if (reset) begin
      ConfReg_10 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_611) begin
              if (_T_642) begin
                if (io_mainMemio_we) begin
                  if (_T_647) begin
                    if (4'ha == confaddr) begin
                      ConfReg_10 <= _T_656;
                    end
                  end else begin
                    if (4'ha == confaddr) begin
                      ConfReg_10 <= _T_644;
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'ha == confaddr) begin
                          ConfReg_10 <= _T_656;
                        end
                      end else begin
                        if (4'ha == confaddr) begin
                          ConfReg_10 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (cond1) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'ha == confaddr) begin
                            ConfReg_10 <= _T_656;
                          end
                        end else begin
                          if (4'ha == confaddr) begin
                            ConfReg_10 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_283) begin
                    if (_T_611) begin
                      if (_T_642) begin
                        if (io_mainMemio_we) begin
                          if (_T_647) begin
                            if (4'ha == confaddr) begin
                              ConfReg_10 <= _T_656;
                            end
                          end else begin
                            if (4'ha == confaddr) begin
                              ConfReg_10 <= _T_644;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        ConfReg_10 <= _T_810;
                      end else begin
                        ConfReg_10 <= _GEN_111;
                      end
                    end else begin
                      ConfReg_10 <= _GEN_111;
                    end
                  end
                end
              end
            end else begin
              ConfReg_10 <= _GEN_111;
            end
          end
        end else begin
          ConfReg_10 <= _GEN_111;
        end
      end else begin
        ConfReg_10 <= _GEN_111;
      end
    end
    if (reset) begin
      ConfReg_11 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_611) begin
              if (_T_642) begin
                if (io_mainMemio_we) begin
                  if (_T_647) begin
                    if (4'hb == confaddr) begin
                      ConfReg_11 <= _T_656;
                    end
                  end else begin
                    if (4'hb == confaddr) begin
                      ConfReg_11 <= _T_644;
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'hb == confaddr) begin
                          ConfReg_11 <= _T_656;
                        end
                      end else begin
                        if (4'hb == confaddr) begin
                          ConfReg_11 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (cond1) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'hb == confaddr) begin
                            ConfReg_11 <= _T_656;
                          end
                        end else begin
                          if (4'hb == confaddr) begin
                            ConfReg_11 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_283) begin
                    if (_T_611) begin
                      if (_T_642) begin
                        if (io_mainMemio_we) begin
                          if (_T_647) begin
                            if (4'hb == confaddr) begin
                              ConfReg_11 <= _T_656;
                            end
                          end else begin
                            if (4'hb == confaddr) begin
                              ConfReg_11 <= _T_644;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        ConfReg_11 <= _T_811;
                      end else begin
                        ConfReg_11 <= _GEN_112;
                      end
                    end else begin
                      ConfReg_11 <= _GEN_112;
                    end
                  end
                end
              end
            end else begin
              ConfReg_11 <= _GEN_112;
            end
          end
        end else begin
          ConfReg_11 <= _GEN_112;
        end
      end else begin
        ConfReg_11 <= _GEN_112;
      end
    end
    if (reset) begin
      ConfReg_12 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_611) begin
              if (_T_642) begin
                if (io_mainMemio_we) begin
                  if (_T_647) begin
                    if (4'hc == confaddr) begin
                      ConfReg_12 <= _T_656;
                    end
                  end else begin
                    if (4'hc == confaddr) begin
                      ConfReg_12 <= _T_644;
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'hc == confaddr) begin
                          ConfReg_12 <= _T_656;
                        end
                      end else begin
                        if (4'hc == confaddr) begin
                          ConfReg_12 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (cond1) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'hc == confaddr) begin
                            ConfReg_12 <= _T_656;
                          end
                        end else begin
                          if (4'hc == confaddr) begin
                            ConfReg_12 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_283) begin
                    if (_T_611) begin
                      if (_T_642) begin
                        if (io_mainMemio_we) begin
                          if (_T_647) begin
                            if (4'hc == confaddr) begin
                              ConfReg_12 <= _T_656;
                            end
                          end else begin
                            if (4'hc == confaddr) begin
                              ConfReg_12 <= _T_644;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        ConfReg_12 <= _T_812;
                      end else begin
                        ConfReg_12 <= _GEN_113;
                      end
                    end else begin
                      ConfReg_12 <= _GEN_113;
                    end
                  end
                end
              end
            end else begin
              ConfReg_12 <= _GEN_113;
            end
          end
        end else begin
          ConfReg_12 <= _GEN_113;
        end
      end else begin
        ConfReg_12 <= _GEN_113;
      end
    end
    if (reset) begin
      ConfReg_13 <= 32'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_611) begin
              if (_T_642) begin
                if (io_mainMemio_we) begin
                  if (_T_647) begin
                    if (4'hd == confaddr) begin
                      ConfReg_13 <= _T_656;
                    end
                  end else begin
                    if (4'hd == confaddr) begin
                      ConfReg_13 <= _T_644;
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_611) begin
                  if (_T_642) begin
                    if (io_mainMemio_we) begin
                      if (_T_647) begin
                        if (4'hd == confaddr) begin
                          ConfReg_13 <= _T_656;
                        end
                      end else begin
                        if (4'hd == confaddr) begin
                          ConfReg_13 <= _T_644;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (cond1) begin
                  if (_T_611) begin
                    if (_T_642) begin
                      if (io_mainMemio_we) begin
                        if (_T_647) begin
                          if (4'hd == confaddr) begin
                            ConfReg_13 <= _T_656;
                          end
                        end else begin
                          if (4'hd == confaddr) begin
                            ConfReg_13 <= _T_644;
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_283) begin
                    if (_T_611) begin
                      if (_T_642) begin
                        if (io_mainMemio_we) begin
                          if (_T_647) begin
                            if (4'hd == confaddr) begin
                              ConfReg_13 <= _T_656;
                            end
                          end else begin
                            if (4'hd == confaddr) begin
                              ConfReg_13 <= _T_644;
                            end
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        ConfReg_13 <= _T_813;
                      end else begin
                        ConfReg_13 <= _GEN_114;
                      end
                    end else begin
                      ConfReg_13 <= _GEN_114;
                    end
                  end
                end
              end
            end else begin
              ConfReg_13 <= _GEN_114;
            end
          end
        end else begin
          ConfReg_13 <= _GEN_114;
        end
      end else begin
        ConfReg_13 <= _GEN_114;
      end
    end
    if (reset) begin
      initState <= 3'h0;
    end else begin
      initState <= initStateNext;
    end
    if (reset) begin
      initStateNext <= 3'h0;
    end else begin
      if (!(moduleReady)) begin
        if (_T_937) begin
          initStateNext <= 3'h1;
        end else begin
          if (_T_938) begin
            if (rndgenm_io_done) begin
              initStateNext <= 3'h2;
            end
          end else begin
            if (_T_939) begin
              if (rndgenm_io_done) begin
                initStateNext <= 3'h3;
              end
            end else begin
              if (_T_940) begin
                if (rndgenm_io_done) begin
                  initStateNext <= 3'h4;
                end
              end else begin
                if (_T_274) begin
                  if (rndgenm_io_done) begin
                    initStateNext <= 3'h5;
                  end
                end else begin
                  if (_T_522) begin
                    if (aesm_io_newR) begin
                      initStateNext <= 3'h6;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      poState <= 3'h6;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (_T_773) begin
              if (_T_342) begin
                poState <= 3'h0;
              end else begin
                if (_T_316) begin
                  poState <= 3'h2;
                end else begin
                  if (_T_359) begin
                    if (aesm_io_newR) begin
                      if (cond2) begin
                        if (_T_253) begin
                          poState <= 3'h1;
                        end else begin
                          poState <= 3'h4;
                        end
                      end else begin
                        poState <= 3'h4;
                      end
                    end else begin
                      poState <= 3'h2;
                    end
                  end else begin
                    if (_T_766) begin
                      if (poutdataReady) begin
                        if (cond2) begin
                          poState <= 3'h1;
                        end else begin
                          poState <= 3'h5;
                        end
                      end else begin
                        poState <= 3'h4;
                      end
                    end else begin
                      if (_T_330) begin
                        if (_T_219) begin
                          if (io_memio_ready) begin
                            poState <= 3'h2;
                          end else begin
                            poState <= 3'h1;
                          end
                        end else begin
                          poState <= 3'h2;
                        end
                      end else begin
                        if (_T_318) begin
                          if (_T_311) begin
                            poState <= 3'h6;
                          end else begin
                            poState <= 3'h5;
                          end
                        end else begin
                          poState <= 3'h6;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              poState <= 3'h6;
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                poState <= 3'h0;
              end else begin
                if (cond1) begin
                  poState <= 3'h1;
                end else begin
                  if (_T_283) begin
                    if (pindataReady) begin
                      poState <= 3'h2;
                    end else begin
                      if (_T_773) begin
                        if (_T_342) begin
                          poState <= 3'h0;
                        end else begin
                          if (_T_316) begin
                            poState <= 3'h2;
                          end else begin
                            if (_T_359) begin
                              if (aesm_io_newR) begin
                                if (cond2) begin
                                  if (_T_253) begin
                                    poState <= 3'h1;
                                  end else begin
                                    poState <= 3'h4;
                                  end
                                end else begin
                                  poState <= 3'h4;
                                end
                              end else begin
                                poState <= 3'h2;
                              end
                            end else begin
                              if (_T_766) begin
                                if (poutdataReady) begin
                                  if (cond2) begin
                                    poState <= 3'h1;
                                  end else begin
                                    poState <= 3'h5;
                                  end
                                end else begin
                                  poState <= 3'h4;
                                end
                              end else begin
                                if (_T_330) begin
                                  if (_T_219) begin
                                    if (io_memio_ready) begin
                                      poState <= 3'h2;
                                    end else begin
                                      poState <= 3'h1;
                                    end
                                  end else begin
                                    poState <= 3'h2;
                                  end
                                end else begin
                                  if (_T_318) begin
                                    if (_T_311) begin
                                      poState <= 3'h6;
                                    end else begin
                                      poState <= 3'h5;
                                    end
                                  end else begin
                                    poState <= 3'h6;
                                  end
                                end
                              end
                            end
                          end
                        end
                      end else begin
                        poState <= 3'h6;
                      end
                    end
                  end else begin
                    if (_T_462) begin
                      if (aesm_io_newR) begin
                        poState <= 3'h3;
                      end else begin
                        if (_T_773) begin
                          if (_T_342) begin
                            poState <= 3'h0;
                          end else begin
                            if (_T_316) begin
                              poState <= 3'h2;
                            end else begin
                              if (_T_359) begin
                                if (aesm_io_newR) begin
                                  if (cond2) begin
                                    if (_T_253) begin
                                      poState <= 3'h1;
                                    end else begin
                                      poState <= 3'h4;
                                    end
                                  end else begin
                                    poState <= 3'h4;
                                  end
                                end else begin
                                  poState <= 3'h2;
                                end
                              end else begin
                                if (_T_766) begin
                                  if (poutdataReady) begin
                                    if (cond2) begin
                                      poState <= 3'h1;
                                    end else begin
                                      poState <= 3'h5;
                                    end
                                  end else begin
                                    poState <= 3'h4;
                                  end
                                end else begin
                                  if (_T_330) begin
                                    if (_T_219) begin
                                      if (io_memio_ready) begin
                                        poState <= 3'h2;
                                      end else begin
                                        poState <= 3'h1;
                                      end
                                    end else begin
                                      poState <= 3'h2;
                                    end
                                  end else begin
                                    if (_T_318) begin
                                      if (_T_311) begin
                                        poState <= 3'h6;
                                      end else begin
                                        poState <= 3'h5;
                                      end
                                    end else begin
                                      poState <= 3'h6;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end else begin
                          poState <= 3'h6;
                        end
                      end
                    end else begin
                      if (_T_436) begin
                        if (_T_894) begin
                          poState <= 3'h2;
                        end else begin
                          if (_T_627) begin
                            if (io_memio_ready) begin
                              if (_T_901) begin
                                poState <= 3'h1;
                              end else begin
                                poState <= 3'h5;
                              end
                            end else begin
                              if (_T_773) begin
                                if (_T_342) begin
                                  poState <= 3'h0;
                                end else begin
                                  if (_T_316) begin
                                    poState <= 3'h2;
                                  end else begin
                                    if (_T_359) begin
                                      if (aesm_io_newR) begin
                                        if (cond2) begin
                                          if (_T_253) begin
                                            poState <= 3'h1;
                                          end else begin
                                            poState <= 3'h4;
                                          end
                                        end else begin
                                          poState <= 3'h4;
                                        end
                                      end else begin
                                        poState <= 3'h2;
                                      end
                                    end else begin
                                      if (_T_766) begin
                                        if (poutdataReady) begin
                                          if (cond2) begin
                                            poState <= 3'h1;
                                          end else begin
                                            poState <= 3'h5;
                                          end
                                        end else begin
                                          poState <= 3'h4;
                                        end
                                      end else begin
                                        if (_T_330) begin
                                          if (_T_219) begin
                                            if (io_memio_ready) begin
                                              poState <= 3'h2;
                                            end else begin
                                              poState <= 3'h1;
                                            end
                                          end else begin
                                            poState <= 3'h2;
                                          end
                                        end else begin
                                          if (_T_318) begin
                                            if (_T_311) begin
                                              poState <= 3'h6;
                                            end else begin
                                              poState <= 3'h5;
                                            end
                                          end else begin
                                            poState <= 3'h6;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end else begin
                                poState <= 3'h6;
                              end
                            end
                          end else begin
                            if (_T_901) begin
                              poState <= 3'h1;
                            end else begin
                              poState <= 3'h5;
                            end
                          end
                        end
                      end else begin
                        if (_T_378) begin
                          if (_T_263) begin
                            poState <= _T_774;
                          end else begin
                            if (_T_835) begin
                              poState <= _T_774;
                            end else begin
                              if (_T_311) begin
                                poState <= 3'h6;
                              end else begin
                                poState <= _T_774;
                              end
                            end
                          end
                        end else begin
                          poState <= _T_774;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              poState <= _T_774;
            end
          end
        end else begin
          poState <= _T_774;
        end
      end else begin
        poState <= _T_774;
      end
    end
    if (reset) begin
      cleanupState <= 2'h0;
    end else begin
      cleanupState <= cleanupStateNext;
    end
    if (reset) begin
      cleanupStateNext <= 2'h0;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (!(_T_290)) begin
              if (cond1) begin
                if (_T_221) begin
                  cleanupStateNext <= 2'h0;
                end
              end else begin
                if (!(_T_283)) begin
                  if (!(_T_462)) begin
                    if (!(_T_823)) begin
                      if (_T_378) begin
                        if (_T_263) begin
                          cleanupStateNext <= 2'h1;
                        end else begin
                          if (_T_835) begin
                            cleanupStateNext <= 2'h2;
                          end else begin
                            if (_T_311) begin
                              cleanupStateNext <= 2'h0;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (_T_290) begin
                if (_T_629) begin
                  cleanupStateNext <= 2'h0;
                end
              end else begin
                if (!(cond1)) begin
                  if (!(_T_283)) begin
                    if (!(_T_462)) begin
                      if (!(_T_436)) begin
                        if (_T_378) begin
                          if (_T_263) begin
                            cleanupStateNext <= 2'h1;
                          end else begin
                            if (_T_835) begin
                              cleanupStateNext <= 2'h2;
                            end else begin
                              if (_T_311) begin
                                cleanupStateNext <= 2'h0;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tagState <= 2'h1;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (!(_T_290)) begin
              if (!(cond1)) begin
                if (_T_283) begin
                  tagState <= 2'h2;
                end else begin
                  if (!(_T_462)) begin
                    if (!(_T_823)) begin
                      if (_T_378) begin
                        if (_T_263) begin
                          tagState <= 2'h3;
                        end else begin
                          if (_T_835) begin
                            tagState <= 2'h1;
                          end else begin
                            if (_T_311) begin
                              tagState <= 2'h1;
                            end else begin
                              tagState <= 2'h3;
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_630) begin
              if (!(_T_290)) begin
                if (!(cond1)) begin
                  if (!(_T_283)) begin
                    if (!(_T_462)) begin
                      if (_T_436) begin
                        tagState <= 2'h2;
                      end else begin
                        if (_T_378) begin
                          if (_T_263) begin
                            tagState <= 2'h3;
                          end else begin
                            if (_T_835) begin
                              tagState <= 2'h1;
                            end else begin
                              if (_T_311) begin
                                tagState <= 2'h1;
                              end else begin
                                tagState <= 2'h3;
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      tagUp <= 1'h1;
    end else begin
      if (moduleReady) begin
        if (start) begin
          if (_T_222) begin
            if (!(_T_290)) begin
              if (!(cond1)) begin
                if (!(_T_283)) begin
                  if (_T_462) begin
                    if (aesm_io_newR) begin
                      tagUp <= 1'h1;
                    end
                  end else begin
                    if (_T_823) begin
                      tagUp <= 1'h0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      encry <= 1'h0;
    end else begin
      if (_T_251) begin
        encry <= _T_522;
      end else begin
        encry <= _T_462;
      end
    end
  end
endmodule
module ModuleTop( // @[:@6110.2]
  input         clock, // @[:@6111.4]
  input         reset, // @[:@6112.4]
  input  [13:0] io_io_addr, // @[:@6113.4]
  input         io_io_valid, // @[:@6113.4]
  input  [31:0] io_io_wdata, // @[:@6113.4]
  input         io_io_we, // @[:@6113.4]
  input         io_io_en, // @[:@6113.4]
  output [31:0] io_io_rdata, // @[:@6113.4]
  output        io_io_ready, // @[:@6113.4]
  output        io_done, // @[:@6113.4]
  output        io_err, // @[:@6113.4]
  output        io_currOutReady // @[:@6113.4]
);
  wire  mem_clock; // @[ModuleTop.scala 27:19:@6115.4]
  wire [10:0] mem_io_blockio_addr; // @[ModuleTop.scala 27:19:@6115.4]
  wire [127:0] mem_io_blockio_wdata; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_blockio_we; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_blockio_en; // @[ModuleTop.scala 27:19:@6115.4]
  wire [127:0] mem_io_blockio_rdata; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_blockio_ready; // @[ModuleTop.scala 27:19:@6115.4]
  wire [12:0] mem_io_dataio_addr; // @[ModuleTop.scala 27:19:@6115.4]
  wire [31:0] mem_io_dataio_wdata; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_dataio_we; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_dataio_en; // @[ModuleTop.scala 27:19:@6115.4]
  wire [31:0] mem_io_dataio_rdata; // @[ModuleTop.scala 27:19:@6115.4]
  wire  mem_io_dataio_ready; // @[ModuleTop.scala 27:19:@6115.4]
  wire  ps_clock; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_reset; // @[ModuleTop.scala 28:19:@6118.4]
  wire [13:0] ps_io_mainMemio_addr; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_mainMemio_valid; // @[ModuleTop.scala 28:19:@6118.4]
  wire [31:0] ps_io_mainMemio_wdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_mainMemio_we; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_mainMemio_en; // @[ModuleTop.scala 28:19:@6118.4]
  wire [31:0] ps_io_mainMemio_rdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_mainMemio_ready; // @[ModuleTop.scala 28:19:@6118.4]
  wire [13:0] ps_io_socMemio_addr; // @[ModuleTop.scala 28:19:@6118.4]
  wire [31:0] ps_io_socMemio_wdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_socMemio_we; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_socMemio_en; // @[ModuleTop.scala 28:19:@6118.4]
  wire [31:0] ps_io_socMemio_rdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_socMemio_ready; // @[ModuleTop.scala 28:19:@6118.4]
  wire [10:0] ps_io_memio_addr; // @[ModuleTop.scala 28:19:@6118.4]
  wire [127:0] ps_io_memio_wdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_memio_we; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_memio_en; // @[ModuleTop.scala 28:19:@6118.4]
  wire [127:0] ps_io_memio_rdata; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_memio_ready; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_err; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_currOutReady; // @[ModuleTop.scala 28:19:@6118.4]
  wire  ps_io_finished; // @[ModuleTop.scala 28:19:@6118.4]
  Memory4 mem ( // @[ModuleTop.scala 27:19:@6115.4]
    .clock(mem_clock),
    .io_blockio_addr(mem_io_blockio_addr),
    .io_blockio_wdata(mem_io_blockio_wdata),
    .io_blockio_we(mem_io_blockio_we),
    .io_blockio_en(mem_io_blockio_en),
    .io_blockio_rdata(mem_io_blockio_rdata),
    .io_blockio_ready(mem_io_blockio_ready),
    .io_dataio_addr(mem_io_dataio_addr),
    .io_dataio_wdata(mem_io_dataio_wdata),
    .io_dataio_we(mem_io_dataio_we),
    .io_dataio_en(mem_io_dataio_en),
    .io_dataio_rdata(mem_io_dataio_rdata),
    .io_dataio_ready(mem_io_dataio_ready)
  );
  pageswappergcm ps ( // @[ModuleTop.scala 28:19:@6118.4]
    .clock(ps_clock),
    .reset(ps_reset),
    .io_mainMemio_addr(ps_io_mainMemio_addr),
    .io_mainMemio_valid(ps_io_mainMemio_valid),
    .io_mainMemio_wdata(ps_io_mainMemio_wdata),
    .io_mainMemio_we(ps_io_mainMemio_we),
    .io_mainMemio_en(ps_io_mainMemio_en),
    .io_mainMemio_rdata(ps_io_mainMemio_rdata),
    .io_mainMemio_ready(ps_io_mainMemio_ready),
    .io_socMemio_addr(ps_io_socMemio_addr),
    .io_socMemio_wdata(ps_io_socMemio_wdata),
    .io_socMemio_we(ps_io_socMemio_we),
    .io_socMemio_en(ps_io_socMemio_en),
    .io_socMemio_rdata(ps_io_socMemio_rdata),
    .io_socMemio_ready(ps_io_socMemio_ready),
    .io_memio_addr(ps_io_memio_addr),
    .io_memio_wdata(ps_io_memio_wdata),
    .io_memio_we(ps_io_memio_we),
    .io_memio_en(ps_io_memio_en),
    .io_memio_rdata(ps_io_memio_rdata),
    .io_memio_ready(ps_io_memio_ready),
    .io_err(ps_io_err),
    .io_currOutReady(ps_io_currOutReady),
    .io_finished(ps_io_finished)
  );
  assign io_io_rdata = ps_io_mainMemio_rdata;
  assign io_io_ready = ps_io_mainMemio_ready;
  assign io_done = ps_io_finished;
  assign io_err = ps_io_err;
  assign io_currOutReady = ps_io_currOutReady;
  assign mem_clock = clock;
  assign mem_io_blockio_addr = ps_io_memio_addr;
  assign mem_io_blockio_wdata = ps_io_memio_wdata;
  assign mem_io_blockio_we = ps_io_memio_we;
  assign mem_io_blockio_en = ps_io_memio_en;
  assign mem_io_dataio_addr = ps_io_socMemio_addr[12:0];
  assign mem_io_dataio_wdata = ps_io_socMemio_wdata;
  assign mem_io_dataio_we = ps_io_socMemio_we;
  assign mem_io_dataio_en = ps_io_socMemio_en;
  assign ps_clock = clock;
  assign ps_reset = reset;
  assign ps_io_mainMemio_addr = io_io_addr;
  assign ps_io_mainMemio_valid = io_io_valid;
  assign ps_io_mainMemio_wdata = io_io_wdata;
  assign ps_io_mainMemio_we = io_io_we;
  assign ps_io_mainMemio_en = io_io_en;
  assign ps_io_socMemio_rdata = mem_io_dataio_rdata;
  assign ps_io_socMemio_ready = mem_io_dataio_ready;
  assign ps_io_memio_rdata = mem_io_blockio_rdata;
  assign ps_io_memio_ready = mem_io_blockio_ready;
endmodule
